************************************************************************
* auCdl Netlist:
* 
* Library Name:  ASKA_DIG2
* Top Cell Name: aska_dig
* View Name:     schematic
* Netlisted on:  Sep  9 14:22:28 2024
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.LDD
*.SCALE METER
.PARAM

*.GLOBAL gnd3i!
+        vdd3i!

*.PIN gnd3i!
*+    vdd3i!

************************************************************************
* Library Name: GATES_JI3V
* Cell Name:    invrji3v
* View Name:    schematic
************************************************************************

.SUBCKT invrji3v in out inh_ground_gnd3i inh_power_vdd3i
*.PININFO in:I out:O inh_ground_gnd3i:B inh_power_vdd3i:B
MMP1 out in inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMN1 out in inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
.ENDS

************************************************************************
* Library Name: GATES_JI3V
* Cell Name:    nand2ji3v
* View Name:    schematic
************************************************************************

.SUBCKT nand2ji3v a b out inh_ground_gnd3i inh_power_vdd3i
*.PININFO a:I b:I out:O inh_ground_gnd3i:B inh_power_vdd3i:B
MMP1 out a inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP2 out b inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMN1 out a net25 inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN2 net25 b inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    AND2JI3VX0
* View Name:    cmos_sch
************************************************************************

.SUBCKT AND2JI3VX0 A B Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xinvr_1 net10 Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=700.00n
Xnand2_1 A B net10 inh_ground_gnd3i inh_power_vdd3i / nand2ji3v GT_PDL=350.00n 
+ GT_PDW=560.00n GT_PUL=300.00n GT_PUW=700.00n
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    DFRRQJI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT DFRRQJI3VX1 C D Q RN inh_ground_gnd3i inh_power_vdd3i
*.PININFO C:I D:I RN:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
MM25 MQIB RN inh_power_vdd3i inh_power_vdd3i PE3I W=720.0n L=300n M=1.0 
+ AD=3.456e-13 AS=3.456e-13 PD=2.4e-06 PS=2.4e-06 NRD=0.375 NRS=0.375
MM24 MQIB CI net227 inh_power_vdd3i PE3I W=960.0n L=300n M=1.0 AD=4.608e-13 
+ AS=4.608e-13 PD=2.88e-06 PS=2.88e-06 NRD=0.28125 NRS=0.28125
MM58 SQIB RN inh_power_vdd3i inh_power_vdd3i PE3I W=720.0n L=300n M=1.0 
+ AD=3.456e-13 AS=3.456e-13 PD=2.4e-06 PS=2.4e-06 NRD=0.375 NRS=0.375
MM56 MQI MQIB inh_power_vdd3i inh_power_vdd3i PE3I W=720.0n L=300n M=1.0 
+ AD=3.456e-13 AS=3.456e-13 PD=2.4e-06 PS=2.4e-06 NRD=0.375 NRS=0.375
MM30 net183 MQI inh_power_vdd3i inh_power_vdd3i PE3I W=1u L=300n M=1.0 
+ AD=4.8e-13 AS=4.8e-13 PD=2.96e-06 PS=2.96e-06 NRD=0.27 NRS=0.27
MM23 net227 D inh_power_vdd3i inh_power_vdd3i PE3I W=960.0n L=300n M=1.0 
+ AD=4.608e-13 AS=4.608e-13 PD=2.88e-06 PS=2.88e-06 NRD=0.28125 NRS=0.28125
MM59 net033 SQIB inh_power_vdd3i inh_power_vdd3i PE3I W=720.0n L=300n M=1.0 
+ AD=3.456e-13 AS=3.456e-13 PD=2.4e-06 PS=2.4e-06 NRD=0.375 NRS=0.375
MM36 net191 net033 inh_power_vdd3i inh_power_vdd3i PE3I W=420.0n L=300n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM35 SQIB CI net191 inh_power_vdd3i PE3I W=420.0n L=300n M=1.0 AD=2.016e-13 
+ AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM34Zf MQIB CIB net187 inh_power_vdd3i PE3I W=420.0n L=300n M=1.0 AD=2.016e-13 
+ AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM33 SQIB CIB net183 inh_power_vdd3i PE3I W=1u L=300n M=1.0 AD=4.8e-13 
+ AS=4.8e-13 PD=2.96e-06 PS=2.96e-06 NRD=0.27 NRS=0.27
MM28 net187 MQI inh_power_vdd3i inh_power_vdd3i PE3I W=420.0n L=300n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
Xinvr_3 SQIB Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.41u
Xinvr_2 CIB CI inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=720.00n
Xinvr_1 C CIB inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=720.00n
MM18 MQIB CIB net165 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM17 MQI MQIB inh_ground_gnd3i inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM15 net165 D net168 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM46 SQIB CI net133 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 AD=2.016e-13 
+ AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM19 MQIB CI net125 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 AD=2.016e-13 
+ AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM51 SQIB CIB net145 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM50 net145 net033 net136 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM49q net033 SQIB inh_ground_gnd3i inh_ground_gnd3i NE3I W=420.0n L=350.0n 
+ M=1.0 AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 
+ NRS=0.642857
MM48 net136 RN inh_ground_gnd3i inh_ground_gnd3i NE3I W=890.0n L=350.0n M=1.0 
+ AD=4.272e-13 AS=4.272e-13 PD=2.74e-06 PS=2.74e-06 NRD=0.303371 NRS=0.303371
MM47 net133 MQI net136 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM44 net168 RN inh_ground_gnd3i inh_ground_gnd3i NE3I W=890.0n L=350.0n M=1.0 
+ AD=4.272e-13 AS=4.272e-13 PD=2.74e-06 PS=2.74e-06 NRD=0.303371 NRS=0.303371
MM61 net125 MQI net168 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
.ENDS

************************************************************************
* Library Name: GATES_JI3V
* Cell Name:    nor2ji3v
* View Name:    schematic
************************************************************************

.SUBCKT nor2ji3v a b out inh_ground_gnd3i inh_power_vdd3i
*.PININFO a:I b:I out:O inh_ground_gnd3i:B inh_power_vdd3i:B
MMP1 out a net32 inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP2 net32 b inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMN1 out b inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN2 out a inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    NO2JI3VX0
* View Name:    cmos_sch
************************************************************************

.SUBCKT NO2JI3VX0 A B Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xnor2_1 A B Q inh_ground_gnd3i inh_power_vdd3i / nor2ji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=850.00n
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    NA2JI3VX0
* View Name:    cmos_sch
************************************************************************

.SUBCKT NA2JI3VX0 A B Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xnand2_1 A B Q inh_ground_gnd3i inh_power_vdd3i / nand2ji3v GT_PDL=350.00n 
+ GT_PDW=560.0n GT_PUL=300.00n GT_PUW=700.00n
.ENDS

************************************************************************
* Library Name: GATES_JI3V
* Cell Name:    o22na2ji3v
* View Name:    schematic
************************************************************************

.SUBCKT o22na2ji3v a b c d out inh_ground_gnd3i inh_power_vdd3i
*.PININFO a:I b:I c:I d:I out:O inh_ground_gnd3i:B inh_power_vdd3i:B
MMN3 net6 c inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN1 out a net6 inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN4 net6 d inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN2 out b net6 inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMP4 net21 d inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP3 out c net21 inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP1 out a net22 inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP2 net22 b inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    ON22JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT ON22JI3VX1 A B C D Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I D:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xo22na2_1 A B C D Q inh_ground_gnd3i inh_power_vdd3i / o22na2ji3v 
+ GT_PUL=300.00n GT_PUW=1.41u GT_PDL=350.00n GT_PDW=890.00n
.ENDS

************************************************************************
* Library Name: GATES_JI3V
* Cell Name:    a2no3ji3v
* View Name:    schematic
************************************************************************

.SUBCKT a2no3ji3v a b c d out inh_ground_gnd3i inh_power_vdd3i
*.PININFO a:I b:I c:I d:I out:O inh_ground_gnd3i:B inh_power_vdd3i:B
MMN4 out d inh_ground_gnd3i inh_ground_gnd3i NE3I W=0.75*GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(0.75*GT_PDW) AS=4.8e-07*(0.75*GT_PDW) 
+ PD=2*(4.8e-07+(0.75*GT_PDW)) PS=2.0*(4.8e-07+(0.75*GT_PDW)) 
+ NRD=2.7e-07/(0.75*GT_PDW) NRS=2.7e-07/(0.75*GT_PDW)
MMN3 out c inh_ground_gnd3i inh_ground_gnd3i NE3I W=0.75*GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(0.75*GT_PDW) AS=4.8e-07*(0.75*GT_PDW) 
+ PD=2*(4.8e-07+(0.75*GT_PDW)) PS=2.0*(4.8e-07+(0.75*GT_PDW)) 
+ NRD=2.7e-07/(0.75*GT_PDW) NRS=2.7e-07/(0.75*GT_PDW)
MMN1 out a net19 inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN2 net19 b inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMP1 net10 a inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP4 out d net22 inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP2 net10 b inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP3 net22 c net10 inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    AN211JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT AN211JI3VX1 A B C D Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I D:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xa2no3_1 A B C D Q inh_ground_gnd3i inh_power_vdd3i / a2no3ji3v GT_PUL=300.00n 
+ GT_PUW=1.41u GT_PDL=350.00n GT_PDW=890.00n
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    INJI3VX0
* View Name:    cmos_sch
************************************************************************

.SUBCKT INJI3VX0 A Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xinvr_1 A Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=940.00n
.ENDS

************************************************************************
* Library Name: GATES_JI3V
* Cell Name:    o2na3ji3v
* View Name:    schematic
************************************************************************

.SUBCKT o2na3ji3v a b c d out inh_ground_gnd3i inh_power_vdd3i
*.PININFO a:I b:I c:I d:I out:O inh_ground_gnd3i:B inh_power_vdd3i:B
MMN2 out b net10 inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN1 out a net10 inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN3 net10 c net25 inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN4 net25 d inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMP4 out d inh_power_vdd3i inh_power_vdd3i PE3I W=0.7*GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(0.7*GT_PUW) AS=4.8e-07*(0.7*GT_PUW) PD=2*(4.8e-07+(0.7*GT_PUW)) 
+ PS=2.0*(4.8e-07+(0.7*GT_PUW)) NRD=2.7e-07/(0.7*GT_PUW) 
+ NRS=2.7e-07/(0.7*GT_PUW)
MMP2 net24 b inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP1 out a net24 inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP3 out c inh_power_vdd3i inh_power_vdd3i PE3I W=0.7*GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(0.7*GT_PUW) AS=4.8e-07*(0.7*GT_PUW) PD=2*(4.8e-07+(0.7*GT_PUW)) 
+ PS=2.0*(4.8e-07+(0.7*GT_PUW)) NRD=2.7e-07/(0.7*GT_PUW) 
+ NRS=2.7e-07/(0.7*GT_PUW)
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    ON211JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT ON211JI3VX1 A B C D Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I D:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xo2na3_1 A B C D Q inh_ground_gnd3i inh_power_vdd3i / o2na3ji3v GT_PUL=300.00n 
+ GT_PUW=1.38u GT_PDL=350.00n GT_PDW=900.0n
.ENDS

************************************************************************
* Library Name: GATES_JI3V
* Cell Name:    a2no2ji3v
* View Name:    schematic
************************************************************************

.SUBCKT a2no2ji3v a b c out inh_ground_gnd3i inh_power_vdd3i
*.PININFO a:I b:I c:I out:O inh_ground_gnd3i:B inh_power_vdd3i:B
MMN2 net41 b inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN1 out a net41 inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN3 out c inh_ground_gnd3i inh_ground_gnd3i NE3I W=0.75*GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(0.75*GT_PDW) AS=4.8e-07*(0.75*GT_PDW) 
+ PD=2*(4.8e-07+(0.75*GT_PDW)) PS=2.0*(4.8e-07+(0.75*GT_PDW)) 
+ NRD=2.7e-07/(0.75*GT_PDW) NRS=2.7e-07/(0.75*GT_PDW)
MMP1 net54 a inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP2 net54 b inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP3 out c net54 inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    AN21JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT AN21JI3VX1 A B C Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xa2no2_1 A B C Q inh_ground_gnd3i inh_power_vdd3i / a2no2ji3v GT_PUL=300.00n 
+ GT_PUW=1.41u GT_PDL=350.00n GT_PDW=890.00n
.ENDS

************************************************************************
* Library Name: GATES_JI3V
* Cell Name:    nand3ji3v
* View Name:    schematic
************************************************************************

.SUBCKT nand3ji3v a b c out inh_ground_gnd3i inh_power_vdd3i
*.PININFO a:I b:I c:I out:O inh_ground_gnd3i:B inh_power_vdd3i:B
MMP1 out a inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP3 out c inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP2 out b inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMN1 out a net37 inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN3 net32 c inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN2 net37 b net32 inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    NA3I1JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT NA3I1JI3VX1 AN B C Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO AN:I B:I C:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xnand3_1 C B net5 Q inh_ground_gnd3i inh_power_vdd3i / nand3ji3v 
+ GT_PDL=350.00n GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.0u
Xinvr_1 AN net5 inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=700.0n
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    NA3JI3VX0
* View Name:    cmos_sch
************************************************************************

.SUBCKT NA3JI3VX0 A B C Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xnand3_1 A B C Q inh_ground_gnd3i inh_power_vdd3i / nand3ji3v GT_PDL=350.00n 
+ GT_PDW=700.00n GT_PUL=300.00n GT_PUW=700.00n
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    NO2I1JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT NO2I1JI3VX1 AN B Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO AN:I B:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xnor2_1 B net12 Q inh_ground_gnd3i inh_power_vdd3i / nor2ji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.41u
Xinvr_1 AN net12 inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=700.0n
.ENDS

************************************************************************
* Library Name: GATES_JI3V
* Cell Name:    nand4ji3v
* View Name:    schematic
************************************************************************

.SUBCKT nand4ji3v a b c out d inh_ground_gnd3i inh_power_vdd3i
*.PININFO a:I b:I c:I d:I out:O inh_ground_gnd3i:B inh_power_vdd3i:B
MMN1 out a net15 inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN3 net16 c net14 inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN2 net15 b net16 inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN4 net14 d inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMP1 out a inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP3 out c inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP2 out b inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP4 out d inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    NA4JI3VX0
* View Name:    cmos_sch
************************************************************************

.SUBCKT NA4JI3VX0 A B C D Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I D:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xnand4_1 A B C Q D inh_ground_gnd3i inh_power_vdd3i / nand4ji3v GT_PUL=300.00n 
+ GT_PUW=700.00n GT_PDL=350.00n GT_PDW=800.0n
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    NA22JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT NA22JI3VX1 A B C Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xnand2_2 net05 C Q inh_ground_gnd3i inh_power_vdd3i / nand2ji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.0u
Xnand2_1 A B net05 inh_ground_gnd3i inh_power_vdd3i / nand2ji3v GT_PDL=350.00n 
+ GT_PDW=560.00n GT_PUL=300.00n GT_PUW=700.0n
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    NA2I1JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT NA2I1JI3VX1 AN B Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO AN:I B:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xinvr_1 AN net4 inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=700.0n
Xnand2_1 B net4 Q inh_ground_gnd3i inh_power_vdd3i / nand2ji3v GT_PDL=350.00n 
+ GT_PDW=890.0n GT_PUL=300.00n GT_PUW=1.0u
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    OR2JI3VX0
* View Name:    cmos_sch
************************************************************************

.SUBCKT OR2JI3VX0 A B Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xinvr_1 net10 Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.000n GT_PUW=700.00n
Xnor2_1 A B net10 inh_ground_gnd3i inh_power_vdd3i / nor2ji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=850.00n
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    BUJI3VX12
* View Name:    cmos_sch
************************************************************************

.SUBCKT BUJI3VX12 A Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xinvr_1 A net9 inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=2.4u GT_PUL=300.00n GT_PUW=5.88u
Xinvr_2 net9 Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=7.2u GT_PUL=300.00n GT_PUW=17.64u
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    AND2JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT AND2JI3VX1 A B Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xinvr_1 net10 Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.41u
Xnand2_1 A B net10 inh_ground_gnd3i inh_power_vdd3i / nand2ji3v GT_PDL=350.00n 
+ GT_PDW=560.00n GT_PUL=300.00n GT_PUW=700.00n
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    BUJI3VX8
* View Name:    cmos_sch
************************************************************************

.SUBCKT BUJI3VX8 A Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xinvr_1 A net9 inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=1.78u GT_PUL=300.00n GT_PUW=4.41u
Xinvr_2 net9 Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=5.34u GT_PUL=300.00n GT_PUW=11.76u
.ENDS

************************************************************************
* Library Name: GATES_JI3V
* Cell Name:    o3na2ji3v
* View Name:    schematic
************************************************************************

.SUBCKT o3na2ji3v a b c d out inh_ground_gnd3i inh_power_vdd3i
*.PININFO a:I b:I c:I d:I out:O inh_ground_gnd3i:B inh_power_vdd3i:B
MMN1 net10 a inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN3 net10 b inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN4 net10 c inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN2 out d net10 inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMP2 out d inh_power_vdd3i inh_power_vdd3i PE3I W=0.6*GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(0.6*GT_PUW) AS=4.8e-07*(0.6*GT_PUW) PD=2*(4.8e-07+(0.6*GT_PUW)) 
+ PS=2.0*(4.8e-07+(0.6*GT_PUW)) NRD=2.7e-07/(0.6*GT_PUW) 
+ NRS=2.7e-07/(0.6*GT_PUW)
MMP1 net20 a inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP4 out c net16 inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP3 net16 b net20 inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    ON31JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT ON31JI3VX1 A B C D Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I D:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xo3na2_1 A B C D Q inh_ground_gnd3i inh_power_vdd3i / o3na2ji3v GT_PUL=300.00n 
+ GT_PUW=1.41u GT_PDL=350.00n GT_PDW=890.00n
.ENDS

************************************************************************
* Library Name: GATES_JI3V
* Cell Name:    a22no2ji3v
* View Name:    schematic
************************************************************************

.SUBCKT a22no2ji3v a b c d out inh_ground_gnd3i inh_power_vdd3i
*.PININFO a:I b:I c:I d:I out:O inh_ground_gnd3i:B inh_power_vdd3i:B
MMN1 out a net21 inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN2 net21 b inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN3 out c net22 inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN4 net22 d inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMP1 net11 a inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP2 net11 b inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP4 out d net11 inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP3 out c net11 inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    AN22JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT AN22JI3VX1 A B C D Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I D:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xa22no2_1 A B C D Q inh_ground_gnd3i inh_power_vdd3i / a22no2ji3v 
+ GT_PUL=300.000n GT_PUW=1.47u GT_PDL=350.00n GT_PDW=890.00n
.ENDS

************************************************************************
* Library Name: GATES_JI3V
* Cell Name:    o2na2ji3v
* View Name:    schematic
************************************************************************

.SUBCKT o2na2ji3v a b c out inh_ground_gnd3i inh_power_vdd3i
*.PININFO a:I b:I c:I out:O inh_ground_gnd3i:B inh_power_vdd3i:B
MMN2 net7 b inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN1 net7 a inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN3 out c net7 inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMP1 out a net17 inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP3 out c inh_power_vdd3i inh_power_vdd3i PE3I W=0.7*GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(0.7*GT_PUW) AS=4.8e-07*(0.7*GT_PUW) PD=2*(4.8e-07+(0.7*GT_PUW)) 
+ PS=2.0*(4.8e-07+(0.7*GT_PUW)) NRD=2.7e-07/(0.7*GT_PUW) 
+ NRS=2.7e-07/(0.7*GT_PUW)
MMP2 net17 b inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    ON21JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT ON21JI3VX1 A B C Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xo2na2_1 A B C Q inh_ground_gnd3i inh_power_vdd3i / o2na2ji3v GT_PUL=300.00n 
+ GT_PUW=1.41u GT_PDL=350.00n GT_PDW=890.00n
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    DFRRQJI3VX4
* View Name:    cmos_sch
************************************************************************

.SUBCKT DFRRQJI3VX4 C D Q RN inh_ground_gnd3i inh_power_vdd3i
*.PININFO C:I D:I RN:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
MM25 MQIB RN inh_power_vdd3i inh_power_vdd3i PE3I W=720.0n L=300n M=1.0 
+ AD=3.456e-13 AS=3.456e-13 PD=2.4e-06 PS=2.4e-06 NRD=0.375 NRS=0.375
MM24 MQIB CI net227 inh_power_vdd3i PE3I W=960.0n L=300n M=1.0 AD=4.608e-13 
+ AS=4.608e-13 PD=2.88e-06 PS=2.88e-06 NRD=0.28125 NRS=0.28125
MM58 SQIB RN inh_power_vdd3i inh_power_vdd3i PE3I W=720.0n L=300n M=1.0 
+ AD=3.456e-13 AS=3.456e-13 PD=2.4e-06 PS=2.4e-06 NRD=0.375 NRS=0.375
MM56 MQI MQIB inh_power_vdd3i inh_power_vdd3i PE3I W=1.41u L=300n M=1.0 
+ AD=6.768e-13 AS=6.768e-13 PD=3.78e-06 PS=3.78e-06 NRD=0.191489 NRS=0.191489
MM30 net183 MQI inh_power_vdd3i inh_power_vdd3i PE3I W=1u L=300n M=1.0 
+ AD=4.8e-13 AS=4.8e-13 PD=2.96e-06 PS=2.96e-06 NRD=0.27 NRS=0.27
MM23 net227 D inh_power_vdd3i inh_power_vdd3i PE3I W=960.0n L=300n M=1.0 
+ AD=4.608e-13 AS=4.608e-13 PD=2.88e-06 PS=2.88e-06 NRD=0.28125 NRS=0.28125
MM59 net033 SQIB inh_power_vdd3i inh_power_vdd3i PE3I W=1.41u L=300n M=1.0 
+ AD=6.768e-13 AS=6.768e-13 PD=3.78e-06 PS=3.78e-06 NRD=0.191489 NRS=0.191489
MM36 net191 net033 inh_power_vdd3i inh_power_vdd3i PE3I W=420.0n L=300n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM35 SQIB CI net191 inh_power_vdd3i PE3I W=420.0n L=300n M=1.0 AD=2.016e-13 
+ AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM34Zf MQIB CIB net187 inh_power_vdd3i PE3I W=420.0n L=300n M=1.0 AD=2.016e-13 
+ AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM33 SQIB CIB net183 inh_power_vdd3i PE3I W=1u L=300n M=1.0 AD=4.8e-13 
+ AS=4.8e-13 PD=2.96e-06 PS=2.96e-06 NRD=0.27 NRS=0.27
MM28 net187 MQI inh_power_vdd3i inh_power_vdd3i PE3I W=420.0n L=300n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
Xinvr_3 SQIB Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=3.56u GT_PUL=300.00n GT_PUW=5.64u
Xinvr_2 CIB CI inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=720.00n
Xinvr_1 C CIB inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=720.00n
MM18 MQIB CIB net165 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM17 MQI MQIB inh_ground_gnd3i inh_ground_gnd3i NE3I W=890.0n L=350.0n M=1.0 
+ AD=4.272e-13 AS=4.272e-13 PD=2.74e-06 PS=2.74e-06 NRD=0.303371 NRS=0.303371
MM15 net165 D net168 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM46 SQIB CI net133 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 AD=2.016e-13 
+ AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM19 MQIB CI net125 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 AD=2.016e-13 
+ AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM51 SQIB CIB net145 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM50 net145 net033 net136 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM49q net033 SQIB inh_ground_gnd3i inh_ground_gnd3i NE3I W=890.0n L=350.0n 
+ M=1.0 AD=4.272e-13 AS=4.272e-13 PD=2.74e-06 PS=2.74e-06 NRD=0.303371 
+ NRS=0.303371
MM48 net136 RN inh_ground_gnd3i inh_ground_gnd3i NE3I W=890.0n L=350.0n M=1.0 
+ AD=4.272e-13 AS=4.272e-13 PD=2.74e-06 PS=2.74e-06 NRD=0.303371 NRS=0.303371
MM47 net133 MQI net136 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM44 net168 RN inh_ground_gnd3i inh_ground_gnd3i NE3I W=890.0n L=350.0n M=1.0 
+ AD=4.272e-13 AS=4.272e-13 PD=2.74e-06 PS=2.74e-06 NRD=0.303371 NRS=0.303371
MM61 net125 MQI net168 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
.ENDS

************************************************************************
* Library Name: GATES_JI3V
* Cell Name:    a2no2_0ji3v
* View Name:    schematic
************************************************************************

.SUBCKT a2no2_0ji3v a b c out inh_ground_gnd3i inh_power_vdd3i
*.PININFO a:I b:I c:I out:O inh_ground_gnd3i:B inh_power_vdd3i:B
MMP1 net54 a inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP2 net54 b inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP3 out c net54 inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMN2 net41 b inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN1 out a net41 inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN3 out c inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    AO21JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT AO21JI3VX1 A B C Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xinvr_1 net15 Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.41u
Xa2no2_1 A B C net15 inh_ground_gnd3i inh_power_vdd3i / a2no2_0ji3v 
+ GT_PDL=350.00n GT_PDW=560.0n GT_PUL=300.00n GT_PUW=850.00n
.ENDS

************************************************************************
* Library Name: GATES_JI3V
* Cell Name:    nor3ji3v
* View Name:    schematic
************************************************************************

.SUBCKT nor3ji3v a b c out inh_ground_gnd3i inh_power_vdd3i
*.PININFO a:I b:I c:I out:O inh_ground_gnd3i:B inh_power_vdd3i:B
MMP3 net37 c inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP1 out a net32 inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP2 net32 b net37 inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMN1 out a inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN3 out c inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN2 out b inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    OR3JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT OR3JI3VX1 A B C Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xinvr_1 net17 Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.41u
Xnor3_1 A B C net17 inh_ground_gnd3i inh_power_vdd3i / nor3ji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=1.00u
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    NO3JI3VX0
* View Name:    cmos_sch
************************************************************************

.SUBCKT NO3JI3VX0 A B C Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xnor3_1 A B C Q inh_ground_gnd3i inh_power_vdd3i / nor3ji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=1.00u
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    NO3I1JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT NO3I1JI3VX1 AN B C Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO AN:I B:I C:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xnor3_1 C B net17 Q inh_ground_gnd3i inh_power_vdd3i / nor3ji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.41u
Xinvr_1 AN net17 inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=700.0n
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    AO22JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT AO22JI3VX1 A B C D Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I D:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xinvr_1 net14 Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.000n GT_PUW=1.47u
Xa22no2_1 A B C D net14 inh_ground_gnd3i inh_power_vdd3i / a22no2ji3v 
+ GT_PUL=300.00n GT_PUW=850.00n GT_PDL=350.00n GT_PDW=560.0n
.ENDS

************************************************************************
* Library Name: GATES_JI3V
* Cell Name:    a3no2ji3v
* View Name:    schematic
************************************************************************

.SUBCKT a3no2ji3v a b c d out inh_ground_gnd3i inh_power_vdd3i
*.PININFO a:I b:I c:I d:I out:O inh_ground_gnd3i:B inh_power_vdd3i:B
MMN3 out c net22 inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN2 out d inh_ground_gnd3i inh_ground_gnd3i NE3I W=0.65*GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(0.65*GT_PDW) AS=4.8e-07*(0.65*GT_PDW) 
+ PD=2*(4.8e-07+(0.65*GT_PDW)) PS=2.0*(4.8e-07+(0.65*GT_PDW)) 
+ NRD=2.7e-07/(0.65*GT_PDW) NRS=2.7e-07/(0.65*GT_PDW)
MMN1 net23 a inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN4 net22 b net23 inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMP3 net10 c inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP4 net10 b inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP1 net10 a inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP2 out d net10 inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    AN31JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT AN31JI3VX1 A B C D Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I D:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xa3no2_1 A B C D Q inh_ground_gnd3i inh_power_vdd3i / a3no2ji3v 
+ GT_PUL=300.000n GT_PUW=1.45u GT_PDL=350.00n GT_PDW=890.0n
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    EO2JI3VX0
* View Name:    cmos_sch
************************************************************************

.SUBCKT EO2JI3VX0 A B Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xnor2_1 A B net10 inh_ground_gnd3i inh_power_vdd3i / nor2ji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=900.00n
Xa2no2_1 A B net10 Q inh_ground_gnd3i inh_power_vdd3i / a2no2_0ji3v 
+ GT_PDL=350.00n GT_PDW=420.00n GT_PUL=300.00n GT_PUW=1.3u
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    FAJI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT FAJI3VX1 A B CI CO S inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I CI:I CO:O S:O inh_ground_gnd3i:B inh_power_vdd3i:B
MM19 net167 CI net99 inh_power_vdd3i PE3I W=1u L=300n M=1.0 AD=4.8e-13 
+ AS=4.8e-13 PD=2.96e-06 PS=2.96e-06 NRD=0.27 NRS=0.27
MM27 net125 A inh_power_vdd3i inh_power_vdd3i PE3I W=1.03u L=300n M=1.0 
+ AD=4.944e-13 AS=4.944e-13 PD=3.02e-06 PS=3.02e-06 NRD=0.262136 NRS=0.262136
MM26 net159 CI net129 inh_power_vdd3i PE3I W=1.03u L=300n M=1.0 AD=4.944e-13 
+ AS=4.944e-13 PD=3.02e-06 PS=3.02e-06 NRD=0.262136 NRS=0.262136
MM25 net129 B net125 inh_power_vdd3i PE3I W=1.03u L=300n M=1.0 AD=4.944e-13 
+ AS=4.944e-13 PD=3.02e-06 PS=3.02e-06 NRD=0.262136 NRS=0.262136
MM24 net159 net167 net107 inh_power_vdd3i PE3I W=1.03u L=300n M=1.0 
+ AD=4.944e-13 AS=4.944e-13 PD=3.02e-06 PS=3.02e-06 NRD=0.262136 NRS=0.262136
MM23 net107 B inh_power_vdd3i inh_power_vdd3i PE3I W=1.03u L=300n M=1.0 
+ AD=4.944e-13 AS=4.944e-13 PD=3.02e-06 PS=3.02e-06 NRD=0.262136 NRS=0.262136
MM22 net107 A inh_power_vdd3i inh_power_vdd3i PE3I W=1.03u L=300n M=1.0 
+ AD=4.944e-13 AS=4.944e-13 PD=3.02e-06 PS=3.02e-06 NRD=0.262136 NRS=0.262136
MM21 net107 CI inh_power_vdd3i inh_power_vdd3i PE3I W=1.03u L=300n M=1.0 
+ AD=4.944e-13 AS=4.944e-13 PD=3.02e-06 PS=3.02e-06 NRD=0.262136 NRS=0.262136
MM20 net99 B inh_power_vdd3i inh_power_vdd3i PE3I W=1u L=300n M=1.0 AD=4.8e-13 
+ AS=4.8e-13 PD=2.96e-06 PS=2.96e-06 NRD=0.27 NRS=0.27
MM18 net99 A inh_power_vdd3i inh_power_vdd3i PE3I W=1u L=300n M=1.0 AD=4.8e-13 
+ AS=4.8e-13 PD=2.96e-06 PS=2.96e-06 NRD=0.27 NRS=0.27
MM17 net167 B net97 inh_power_vdd3i PE3I W=1u L=300n M=1.0 AD=4.8e-13 
+ AS=4.8e-13 PD=2.96e-06 PS=2.96e-06 NRD=0.27 NRS=0.27
MM16 net97 A inh_power_vdd3i inh_power_vdd3i PE3I W=1u L=300n M=1.0 AD=4.8e-13 
+ AS=4.8e-13 PD=2.96e-06 PS=2.96e-06 NRD=0.27 NRS=0.27
MM8 net175 A inh_ground_gnd3i inh_ground_gnd3i NE3I W=550.0n L=350.0n M=1.0 
+ AD=2.64e-13 AS=2.64e-13 PD=2.06e-06 PS=2.06e-06 NRD=0.490909 NRS=0.490909
MM10 net179 A inh_ground_gnd3i inh_ground_gnd3i NE3I W=590.0n L=350.0n M=1.0 
+ AD=2.832e-13 AS=2.832e-13 PD=2.14e-06 PS=2.14e-06 NRD=0.457627 NRS=0.457627
MM6 net175 CI inh_ground_gnd3i inh_ground_gnd3i NE3I W=550.0n L=350.0n M=1.0 
+ AD=2.64e-13 AS=2.64e-13 PD=2.06e-06 PS=2.06e-06 NRD=0.490909 NRS=0.490909
MM11 net171 B net179 inh_ground_gnd3i NE3I W=590.0n L=350.0n M=1.0 
+ AD=2.832e-13 AS=2.832e-13 PD=2.14e-06 PS=2.14e-06 NRD=0.457627 NRS=0.457627
MM1 net167 B net151 inh_ground_gnd3i NE3I W=590.0n L=350.0n M=1.0 AD=2.832e-13 
+ AS=2.832e-13 PD=2.14e-06 PS=2.14e-06 NRD=0.457627 NRS=0.457627
MM4 net163 A inh_ground_gnd3i inh_ground_gnd3i NE3I W=590.0n L=350.0n M=1.0 
+ AD=2.832e-13 AS=2.832e-13 PD=2.14e-06 PS=2.14e-06 NRD=0.457627 NRS=0.457627
MM9 net159 net167 net175 inh_ground_gnd3i NE3I W=480.0n L=350.0n M=1.0 
+ AD=2.304e-13 AS=2.304e-13 PD=1.92e-06 PS=1.92e-06 NRD=0.5625 NRS=0.5625
MM3 net167 CI net163 inh_ground_gnd3i NE3I W=590.0n L=350.0n M=1.0 
+ AD=2.832e-13 AS=2.832e-13 PD=2.14e-06 PS=2.14e-06 NRD=0.457627 NRS=0.457627
MM2 net151 A inh_ground_gnd3i inh_ground_gnd3i NE3I W=590.0n L=350.0n M=1.0 
+ AD=2.832e-13 AS=2.832e-13 PD=2.14e-06 PS=2.14e-06 NRD=0.457627 NRS=0.457627
MM12 net159 CI net171 inh_ground_gnd3i NE3I W=590.0n L=350.0n M=1.0 
+ AD=2.832e-13 AS=2.832e-13 PD=2.14e-06 PS=2.14e-06 NRD=0.457627 NRS=0.457627
MM7 net175 B inh_ground_gnd3i inh_ground_gnd3i NE3I W=480.0n L=350.0n M=1.0 
+ AD=2.304e-13 AS=2.304e-13 PD=1.92e-06 PS=1.92e-06 NRD=0.5625 NRS=0.5625
MM5 net163 B inh_ground_gnd3i inh_ground_gnd3i NE3I W=590.0n L=350.0n M=1.0 
+ AD=2.832e-13 AS=2.832e-13 PD=2.14e-06 PS=2.14e-06 NRD=0.457627 NRS=0.457627
Xinvr_2 net159 S inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.41u
Xinvr_1 net167 CO inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=590.00n GT_PUL=300.00n GT_PUW=1.11u
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    BUJI3VX0
* View Name:    cmos_sch
************************************************************************

.SUBCKT BUJI3VX0 A Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xinvr_1 A net9 inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=900.0n
Xinvr_2 net9 Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=1.12u
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    EN3JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT EN3JI3VX1 A B C Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xa2no2_1 B C net19 net29 inh_ground_gnd3i inh_power_vdd3i / a2no2_0ji3v 
+ GT_PDL=350.00n GT_PDW=520.00n GT_PUL=300.00n GT_PUW=1.41u
Xnor2_1 B C net19 inh_ground_gnd3i inh_power_vdd3i / nor2ji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=1.41u
Xo2na2_1 net29 A net16 Q inh_ground_gnd3i inh_power_vdd3i / o2na2ji3v 
+ GT_PUL=300.00n GT_PUW=1.41u GT_PDL=350.00n GT_PDW=420.00n
Xnand2_1 net29 A net16 inh_ground_gnd3i inh_power_vdd3i / nand2ji3v 
+ GT_PDL=350.00n GT_PDW=420.00n GT_PUL=300.00n GT_PUW=1.41u
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    NO3I2JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT NO3I2JI3VX1 AN BN C Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO AN:I BN:I C:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xnand2_1 AN BN net7 inh_ground_gnd3i inh_power_vdd3i / nand2ji3v 
+ GT_PDL=350.00n GT_PDW=480.0n GT_PUL=300.00n GT_PUW=700.0n
Xnor2_1 net7 C Q inh_ground_gnd3i inh_power_vdd3i / nor2ji3v GT_PDL=350.00n 
+ GT_PDW=890.0n GT_PUL=300.00n GT_PUW=1.41u
.ENDS

************************************************************************
* Library Name: GATES_JI3V
* Cell Name:    o2na2_0ji3v
* View Name:    schematic
************************************************************************

.SUBCKT o2na2_0ji3v a b c out inh_ground_gnd3i inh_power_vdd3i
*.PININFO a:I b:I c:I out:O inh_ground_gnd3i:B inh_power_vdd3i:B
MMN2 net7 b inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN1 net7 a inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN3 out c net7 inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMP1 out a net17 inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP3 out c inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP2 net17 b inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    OA21JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT OA21JI3VX1 A B C Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xinvr_1 net15 Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.41u
Xo2na2_1 A B C net15 inh_ground_gnd3i inh_power_vdd3i / o2na2_0ji3v 
+ GT_PUL=300.00n GT_PUW=850.0n GT_PDL=350.00n GT_PDW=540.00n
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    HAJI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT HAJI3VX1 A B CO S inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I CO:O S:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xinvr_2 net49 S inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.41u
Xinvr_1 net64 CO inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=550.00n GT_PUL=300.00n GT_PUW=1.11u
Mmp1 net49 net64 inh_power_vdd3i inh_power_vdd3i PE3I W=890.0n L=300n M=1.0 
+ AD=4.272e-13 AS=4.272e-13 PD=2.74e-06 PS=2.74e-06 NRD=0.303371 NRS=0.303371
Mmp2 net49 B net41 inh_power_vdd3i PE3I W=890.0n L=300n M=1.0 AD=4.272e-13 
+ AS=4.272e-13 PD=2.74e-06 PS=2.74e-06 NRD=0.303371 NRS=0.303371
Mmp3 net41 A inh_power_vdd3i inh_power_vdd3i PE3I W=890.0n L=300n M=1.0 
+ AD=4.272e-13 AS=4.272e-13 PD=2.74e-06 PS=2.74e-06 NRD=0.303371 NRS=0.303371
Xnand2_1 A B net64 inh_ground_gnd3i inh_power_vdd3i / nand2ji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.11u
Mmn3 net53 B inh_ground_gnd3i inh_ground_gnd3i NE3I W=890.0n L=350.0n M=1.0 
+ AD=4.272e-13 AS=4.272e-13 PD=2.74e-06 PS=2.74e-06 NRD=0.303371 NRS=0.303371
Mmn2 net53 A inh_ground_gnd3i inh_ground_gnd3i NE3I W=890.0n L=350.0n M=1.0 
+ AD=4.272e-13 AS=4.272e-13 PD=2.74e-06 PS=2.74e-06 NRD=0.303371 NRS=0.303371
Mmn1 net49 net64 net53 inh_ground_gnd3i NE3I W=590.0n L=350.0n M=1.0 
+ AD=2.832e-13 AS=2.832e-13 PD=2.14e-06 PS=2.14e-06 NRD=0.457627 NRS=0.457627
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    DLY1JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT DLY1JI3VX1 A Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
MM3 net35 net31 inh_power_vdd3i inh_power_vdd3i PE3I W=420.0n L=750.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM1 net31 net47 inh_power_vdd3i inh_power_vdd3i PE3I W=420.0n L=1u M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
Xinvr_2 net35 Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.41u
Xinvr_1 A net47 inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=670.00n
MM2 net31 net47 inh_ground_gnd3i inh_ground_gnd3i NE3I W=420.0n L=800n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM4 net35 net31 inh_ground_gnd3i inh_ground_gnd3i NE3I W=420.0n L=1u M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    NA3I2JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT NA3I2JI3VX1 AN BN C Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO AN:I BN:I C:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xnand2_1 net7 C Q inh_ground_gnd3i inh_power_vdd3i / nand2ji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.0u
Xnor2_1 AN BN net7 inh_ground_gnd3i inh_power_vdd3i / nor2ji3v GT_PDL=350.00n 
+ GT_PDW=420.0n GT_PUL=300.00n GT_PUW=850.00n
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    NO22JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT NO22JI3VX1 A B C Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xnor2_2 net05 C Q inh_ground_gnd3i inh_power_vdd3i / nor2ji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.41u
Xnor2_1 A B net05 inh_ground_gnd3i inh_power_vdd3i / nor2ji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=850.00n
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    EN2JI3VX0
* View Name:    cmos_sch
************************************************************************

.SUBCKT EN2JI3VX0 A B Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xnand2_1 A B net4 inh_ground_gnd3i inh_power_vdd3i / nand2ji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=900.00n
Xo2na2_1 B A net4 Q inh_ground_gnd3i inh_power_vdd3i / o2na2ji3v 
+ GT_PUL=300.00n GT_PUW=1.3u GT_PDL=350.00n GT_PDW=420.00n
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    SDFRRQJI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT SDFRRQJI3VX1 C D Q RN SD SE inh_ground_gnd3i inh_power_vdd3i
*.PININFO C:I D:I RN:I SD:I SE:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
MM3 MQIB CI net046 inh_power_vdd3i PE3I W=850.0n L=300n M=1.0 AD=4.08e-13 
+ AS=4.08e-13 PD=2.66e-06 PS=2.66e-06 NRD=0.317647 NRS=0.317647
MM22 net061 SE inh_power_vdd3i inh_power_vdd3i PE3I W=900n L=300n M=1.0 
+ AD=4.32e-13 AS=4.32e-13 PD=2.76e-06 PS=2.76e-06 NRD=0.3 NRS=0.3
MM2 net046 D net061 inh_power_vdd3i PE3I W=900n L=300n M=1.0 AD=4.32e-13 
+ AS=4.32e-13 PD=2.76e-06 PS=2.76e-06 NRD=0.3 NRS=0.3
MM26 net046 SD net063 inh_power_vdd3i PE3I W=900n L=300n M=1.0 AD=4.32e-13 
+ AS=4.32e-13 PD=2.76e-06 PS=2.76e-06 NRD=0.3 NRS=0.3
MM21 net063 SEB inh_power_vdd3i inh_power_vdd3i PE3I W=900n L=300n M=1.0 
+ AD=4.32e-13 AS=4.32e-13 PD=2.76e-06 PS=2.76e-06 NRD=0.3 NRS=0.3
MM25 MQIB RN inh_power_vdd3i inh_power_vdd3i PE3I W=1.02u L=300n M=1.0 
+ AD=4.896e-13 AS=4.896e-13 PD=3e-06 PS=3e-06 NRD=0.264706 NRS=0.264706
MM58 SQIB RN inh_power_vdd3i inh_power_vdd3i PE3I W=790.0n L=300n M=1.0 
+ AD=3.792e-13 AS=3.792e-13 PD=2.54e-06 PS=2.54e-06 NRD=0.341772 NRS=0.341772
MM56 MQI MQIB inh_power_vdd3i inh_power_vdd3i PE3I W=1.07u L=300n M=1.0 
+ AD=5.136e-13 AS=5.136e-13 PD=3.1e-06 PS=3.1e-06 NRD=0.252336 NRS=0.252336
MM30 net183 MQI inh_power_vdd3i inh_power_vdd3i PE3I W=790.0n L=300n M=1.0 
+ AD=3.792e-13 AS=3.792e-13 PD=2.54e-06 PS=2.54e-06 NRD=0.341772 NRS=0.341772
MM59 net033 SQIB inh_power_vdd3i inh_power_vdd3i PE3I W=1.41u L=300n M=1.0 
+ AD=6.768e-13 AS=6.768e-13 PD=3.78e-06 PS=3.78e-06 NRD=0.191489 NRS=0.191489
MM36 net191 net033 inh_power_vdd3i inh_power_vdd3i PE3I W=420.0n L=300n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM35 SQIB CI net191 inh_power_vdd3i PE3I W=420.0n L=300n M=1.0 AD=2.016e-13 
+ AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM34 MQIB CIB net187 inh_power_vdd3i PE3I W=420.0n L=300n M=1.0 AD=2.016e-13 
+ AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM33 SQIB CIB net183 inh_power_vdd3i PE3I W=790.0n L=300n M=1.0 AD=3.792e-13 
+ AS=3.792e-13 PD=2.54e-06 PS=2.54e-06 NRD=0.341772 NRS=0.341772
MM28 net187 MQI inh_power_vdd3i inh_power_vdd3i PE3I W=420.0n L=300n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
Xinvr_3 CIB CI inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=720.00n
Xinvr_1 C CIB inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=720.00n
Xinvr_2 SE SEB inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=720.00n
Xinvr_4 SQIB Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.41u
MM1 MQIB CIB net045 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 AD=2.016e-13 
+ AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM16 net062 SEB net168 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM0 net045 D net062 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 AD=2.016e-13 
+ AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM14 net064 SE net168 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM4 net168 RN inh_ground_gnd3i inh_ground_gnd3i NE3I W=540.0n L=350.0n M=1.0 
+ AD=2.592e-13 AS=2.592e-13 PD=2.04e-06 PS=2.04e-06 NRD=0.5 NRS=0.5
MM169 net045 SD net064 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM17 MQI MQIB inh_ground_gnd3i inh_ground_gnd3i NE3I W=720.0n L=350.0n M=1.0 
+ AD=3.456e-13 AS=3.456e-13 PD=2.4e-06 PS=2.4e-06 NRD=0.375 NRS=0.375
MM46 SQIB CI net133 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 AD=2.016e-13 
+ AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM19 MQIB CI net125 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 AD=2.016e-13 
+ AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM51 SQIB CIB net145 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM50 net145 net033 net136 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM49 net033 SQIB inh_ground_gnd3i inh_ground_gnd3i NE3I W=890.0n L=350.0n 
+ M=1.0 AD=4.272e-13 AS=4.272e-13 PD=2.74e-06 PS=2.74e-06 NRD=0.303371 
+ NRS=0.303371
MM48 net136 RN inh_ground_gnd3i inh_ground_gnd3i NE3I W=890.0n L=350.0n M=1.0 
+ AD=4.272e-13 AS=4.272e-13 PD=2.74e-06 PS=2.74e-06 NRD=0.303371 NRS=0.303371
MM47 net133 MQI net136 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM44 net068 RN inh_ground_gnd3i inh_ground_gnd3i NE3I W=890.0n L=350.0n M=1.0 
+ AD=4.272e-13 AS=4.272e-13 PD=2.74e-06 PS=2.74e-06 NRD=0.303371 NRS=0.303371
MM61 net125 MQI net068 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    INJI3VX3
* View Name:    cmos_sch
************************************************************************

.SUBCKT INJI3VX3 A Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xinvr_1 A Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=1.78u GT_PUL=300.00n GT_PUW=4.41u
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    NA4JI3VX2
* View Name:    cmos_sch
************************************************************************

.SUBCKT NA4JI3VX2 A B C D Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I D:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xnand4_1<0> A B C Q D inh_ground_gnd3i inh_power_vdd3i / nand4ji3v 
+ GT_PUL=300.00n GT_PUW=1.00u GT_PDL=350.00n GT_PDW=890.00n
Xnand4_1<1> A B C Q D inh_ground_gnd3i inh_power_vdd3i / nand4ji3v 
+ GT_PUL=300.00n GT_PUW=1.00u GT_PDL=350.00n GT_PDW=890.00n
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    NO2I1JI3VX2
* View Name:    cmos_sch
************************************************************************

.SUBCKT NO2I1JI3VX2 AN B Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO AN:I B:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xnor2_1<0> B net12 Q inh_ground_gnd3i inh_power_vdd3i / nor2ji3v 
+ GT_PDL=350.00n GT_PDW=900.00n GT_PUL=300.00n GT_PUW=1.41u
Xnor2_1<1> B net12 Q inh_ground_gnd3i inh_power_vdd3i / nor2ji3v 
+ GT_PDL=350.00n GT_PDW=900.00n GT_PUL=300.00n GT_PUW=1.41u
Xinvr_1 AN net12 inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=900.00n GT_PUL=300.00n GT_PUW=1.41u
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    OR4JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT OR4JI3VX1 A B C D Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I D:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xnor2_1 C D net21 inh_ground_gnd3i inh_power_vdd3i / nor2ji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=850.0n
Xnor2_2 A B net20 inh_ground_gnd3i inh_power_vdd3i / nor2ji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=850.0n
Xnand2_1 net20 net21 Q inh_ground_gnd3i inh_power_vdd3i / nand2ji3v 
+ GT_PDL=350.00n GT_PDW=890.0n GT_PUL=300.00n GT_PUW=1.41u
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    BUJI3VX2
* View Name:    cmos_sch
************************************************************************

.SUBCKT BUJI3VX2 A Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xinvr_1 A net9 inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=600.00n GT_PUL=300.00n GT_PUW=1.1u
Xinvr_2 net9 Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=1.2u GT_PUL=300.00n GT_PUW=2.92u
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    BUJI3VX3
* View Name:    cmos_sch
************************************************************************

.SUBCKT BUJI3VX3 A Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xinvr_1 A net9 inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.46u
Xinvr_2 net9 Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=1.78u GT_PUL=300.00n GT_PUW=4.38u
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    ON21JI3VX4
* View Name:    cmos_sch
************************************************************************

.SUBCKT ON21JI3VX4 A B C Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xinvr_2<0> net6 Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.43u
Xinvr_2<1> net6 Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.43u
Xinvr_2<2> net6 Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.43u
Xinvr_2<3> net6 Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.43u
Xinvr_1 net5 net6 inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.41u
Xo2na2_1 A B C net5 inh_ground_gnd3i inh_power_vdd3i / o2na2_0ji3v 
+ GT_PUL=300.00n GT_PUW=1.41u GT_PDL=350.00n GT_PDW=890.00n
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    BUJI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT BUJI3VX1 A Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xinvr_1 A net9 inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=900.0n
Xinvr_2 net9 Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=660.0n GT_PUL=300.00n GT_PUW=1.46u
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    INJI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT INJI3VX1 A Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xinvr_1 A Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=600.00n GT_PUL=300.00n GT_PUW=1.41u
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    INJI3VX2
* View Name:    cmos_sch
************************************************************************

.SUBCKT INJI3VX2 A Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xinvr_1 A Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=960.00n GT_PUL=300.00n GT_PUW=2.94u
.ENDS

************************************************************************
* Library Name: GATES_JI3V
* Cell Name:    clinvrji3v
* View Name:    schematic
************************************************************************

.SUBCKT clinvrji3v clk in out xclk inh_ground_gnd3i inh_power_vdd3i
*.PININFO clk:I in:I xclk:I out:O inh_ground_gnd3i:B inh_power_vdd3i:B
MMP2 out xclk net34 inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMP1 net34 in inh_power_vdd3i inh_power_vdd3i PE3I W=GT_PUW L=GT_PUL M=1.0 
+ AD=4.8e-07*(GT_PUW) AS=4.8e-07*(GT_PUW) PD=2*(4.8e-07+(GT_PUW)) 
+ PS=2.0*(4.8e-07+(GT_PUW)) NRD=2.7e-07/(GT_PUW) NRS=2.7e-07/(GT_PUW)
MMN1 net26 in inh_ground_gnd3i inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
MMN2 out clk net26 inh_ground_gnd3i NE3I W=GT_PDW L=GT_PDL M=1.0 
+ AD=4.8e-07*(GT_PDW) AS=4.8e-07*(GT_PDW) PD=2*(4.8e-07+(GT_PDW)) 
+ PS=2.0*(4.8e-07+(GT_PDW)) NRD=2.7e-07/(GT_PDW) NRS=2.7e-07/(GT_PDW)
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    MU2JI3VX0
* View Name:    cmos_sch
************************************************************************

.SUBCKT MU2JI3VX0 IN0 IN1 Q S inh_ground_gnd3i inh_power_vdd3i
*.PININFO IN0:I IN1:I S:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xclinvr_1 S IN1 net22 net20 inh_ground_gnd3i inh_power_vdd3i / clinvrji3v 
+ GT_PDL=350.00n GT_PDW=420.00n GT_PUL=300.00n GT_PUW=780.00n
Xclinvr_2 net20 IN0 net22 S inh_ground_gnd3i inh_power_vdd3i / clinvrji3v 
+ GT_PDL=350.00n GT_PDW=420.00n GT_PUL=300.00n GT_PUW=780.00n
Xinvr_1 S net20 inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=500.00n
Xinvr_2 net22 Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=700.00n
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    BUJI3VX6
* View Name:    cmos_sch
************************************************************************

.SUBCKT BUJI3VX6 A Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xinvr_1 A net9 inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=1.6u GT_PUL=300.00n GT_PUW=2.92u
Xinvr_2 net9 Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=3.56u GT_PUL=300.00n GT_PUW=8.76u
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    NO3JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT NO3JI3VX1 A B C Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xnor3_1 A B C Q inh_ground_gnd3i inh_power_vdd3i / nor3ji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.41u
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    OR4JI3VX2
* View Name:    cmos_sch
************************************************************************

.SUBCKT OR4JI3VX2 A B C D Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I D:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xnor2_1 C D net21 inh_ground_gnd3i inh_power_vdd3i / nor2ji3v GT_PDL=350.00n 
+ GT_PDW=700.00n GT_PUL=300.00n GT_PUW=1.41u
Xnor2_2 A B net20 inh_ground_gnd3i inh_power_vdd3i / nor2ji3v GT_PDL=350.00n 
+ GT_PDW=700.00n GT_PUL=300.00n GT_PUW=1.41u
Xnand2_1<0> net20 net21 Q inh_ground_gnd3i inh_power_vdd3i / nand2ji3v 
+ GT_PDL=350.00n GT_PDW=890.0n GT_PUL=300.00n GT_PUW=1.42u
Xnand2_1<1> net20 net21 Q inh_ground_gnd3i inh_power_vdd3i / nand2ji3v 
+ GT_PDL=350.00n GT_PDW=890.0n GT_PUL=300.00n GT_PUW=1.42u
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    EO3JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT EO3JI3VX1 A B C Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I C:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xa2no2_2 net34 A net24 Q inh_ground_gnd3i inh_power_vdd3i / a2no2_0ji3v 
+ GT_PDL=350.00n GT_PDW=520.00n GT_PUL=300.00n GT_PUW=1.41u
Xa2no2_1 B C net21 net34 inh_ground_gnd3i inh_power_vdd3i / a2no2_0ji3v 
+ GT_PDL=350.00n GT_PDW=520.00n GT_PUL=300.00n GT_PUW=1.41u
Xnor2_1 B C net21 inh_ground_gnd3i inh_power_vdd3i / nor2ji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=1.3u
Xnor2_2 A net34 net24 inh_ground_gnd3i inh_power_vdd3i / nor2ji3v 
+ GT_PDL=350.00n GT_PDW=420.00n GT_PUL=300.00n GT_PUW=1.3u
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    BUJI3VX16
* View Name:    cmos_sch
************************************************************************

.SUBCKT BUJI3VX16 A Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xinvr_1 A net9 inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=4.45u GT_PUL=300.00n GT_PUW=8.82u
Xinvr_2 net9 Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=9.78u GT_PUL=300.00n GT_PUW=23.52u
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    DLY4JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT DLY4JI3VX1 A Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
MM3 net039 net47 net086 inh_power_vdd3i PE3I W=420.0n L=1.2u M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM7 net082 net039 inh_power_vdd3i inh_power_vdd3i PE3I W=420.0n L=1.9u M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM2 net086 net47 inh_power_vdd3i inh_power_vdd3i PE3I W=420.0n L=1.2u M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM8 net35 net039 net082 inh_power_vdd3i PE3I W=420.0n L=1.9u M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
Xinvr_2 net35 Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.41u
Xinvr_1 A net47 inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=700.00n
MM10 net051 net039 inh_ground_gnd3i inh_ground_gnd3i NE3I W=420.0n L=1.1u 
+ M=1.0 AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 
+ NRS=0.642857
MM5 net055 net47 inh_ground_gnd3i inh_ground_gnd3i NE3I W=420.0n L=1.8u M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM9 net35 net039 net051 inh_ground_gnd3i NE3I W=420.0n L=1.1u M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM4 net039 net47 net055 inh_ground_gnd3i NE3I W=420.0n L=1.8u M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    DFRRQJI3VX2
* View Name:    cmos_sch
************************************************************************

.SUBCKT DFRRQJI3VX2 C D Q RN inh_ground_gnd3i inh_power_vdd3i
*.PININFO C:I D:I RN:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
MM25 MQIB RN inh_power_vdd3i inh_power_vdd3i PE3I W=720.0n L=300n M=1.0 
+ AD=3.456e-13 AS=3.456e-13 PD=2.4e-06 PS=2.4e-06 NRD=0.375 NRS=0.375
MM24 MQIB CI net227 inh_power_vdd3i PE3I W=960.0n L=300n M=1.0 AD=4.608e-13 
+ AS=4.608e-13 PD=2.88e-06 PS=2.88e-06 NRD=0.28125 NRS=0.28125
MM58 SQIB RN inh_power_vdd3i inh_power_vdd3i PE3I W=720.0n L=300n M=1.0 
+ AD=3.456e-13 AS=3.456e-13 PD=2.4e-06 PS=2.4e-06 NRD=0.375 NRS=0.375
MM56 MQI MQIB inh_power_vdd3i inh_power_vdd3i PE3I W=1u L=300n M=1.0 
+ AD=4.8e-13 AS=4.8e-13 PD=2.96e-06 PS=2.96e-06 NRD=0.27 NRS=0.27
MM30 net183 MQI inh_power_vdd3i inh_power_vdd3i PE3I W=1u L=300n M=1.0 
+ AD=4.8e-13 AS=4.8e-13 PD=2.96e-06 PS=2.96e-06 NRD=0.27 NRS=0.27
MM23 net227 D inh_power_vdd3i inh_power_vdd3i PE3I W=960.0n L=300n M=1.0 
+ AD=4.608e-13 AS=4.608e-13 PD=2.88e-06 PS=2.88e-06 NRD=0.28125 NRS=0.28125
MM59 net033 SQIB inh_power_vdd3i inh_power_vdd3i PE3I W=1u L=300n M=1.0 
+ AD=4.8e-13 AS=4.8e-13 PD=2.96e-06 PS=2.96e-06 NRD=0.27 NRS=0.27
MM36 net191 net033 inh_power_vdd3i inh_power_vdd3i PE3I W=420.0n L=300n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM35 SQIB CI net191 inh_power_vdd3i PE3I W=420.0n L=300n M=1.0 AD=2.016e-13 
+ AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM34Zf MQIB CIB net187 inh_power_vdd3i PE3I W=420.0n L=300n M=1.0 AD=2.016e-13 
+ AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM33 SQIB CIB net183 inh_power_vdd3i PE3I W=1u L=300n M=1.0 AD=4.8e-13 
+ AS=4.8e-13 PD=2.96e-06 PS=2.96e-06 NRD=0.27 NRS=0.27
MM28 net187 MQI inh_power_vdd3i inh_power_vdd3i PE3I W=420.0n L=300n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
Xinvr_3 SQIB Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=1.78u GT_PUL=300.00n GT_PUW=2.82u
Xinvr_2 CIB CI inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=720.00n
Xinvr_1 C CIB inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=720.00n
MM18 MQIB CIB net165 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM17 MQI MQIB inh_ground_gnd3i inh_ground_gnd3i NE3I W=660.0n L=350.0n M=1.0 
+ AD=3.168e-13 AS=3.168e-13 PD=2.28e-06 PS=2.28e-06 NRD=0.409091 NRS=0.409091
MM15 net165 D net168 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM46 SQIB CI net133 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 AD=2.016e-13 
+ AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM19 MQIB CI net125 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 AD=2.016e-13 
+ AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM51 SQIB CIB net145 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM50 net145 net033 net136 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM49q net033 SQIB inh_ground_gnd3i inh_ground_gnd3i NE3I W=660.0n L=350.0n 
+ M=1.0 AD=3.168e-13 AS=3.168e-13 PD=2.28e-06 PS=2.28e-06 NRD=0.409091 
+ NRS=0.409091
MM48 net136 RN inh_ground_gnd3i inh_ground_gnd3i NE3I W=890.0n L=350.0n M=1.0 
+ AD=4.272e-13 AS=4.272e-13 PD=2.74e-06 PS=2.74e-06 NRD=0.303371 NRS=0.303371
MM47 net133 MQI net136 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM44 net168 RN inh_ground_gnd3i inh_ground_gnd3i NE3I W=890.0n L=350.0n M=1.0 
+ AD=4.272e-13 AS=4.272e-13 PD=2.74e-06 PS=2.74e-06 NRD=0.303371 NRS=0.303371
MM61 net125 MQI net168 inh_ground_gnd3i NE3I W=420.0n L=350.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    DLY2JI3VX1
* View Name:    cmos_sch
************************************************************************

.SUBCKT DLY2JI3VX1 A Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
MM5 net080 net039 inh_power_vdd3i inh_power_vdd3i PE3I W=420.0n L=1u M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM2 net039 net47 net084 inh_power_vdd3i PE3I W=420.0n L=740.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM6 net35 net039 net080 inh_power_vdd3i PE3I W=420.0n L=1u M=1.0 AD=2.016e-13 
+ AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM1 net084 net47 inh_power_vdd3i inh_power_vdd3i PE3I W=420.0n L=740.0n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
Xinvr_2 net35 Q inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.41u
Xinvr_1 A net47 inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=420.00n GT_PUL=300.00n GT_PUW=700.00n
MM4 net31 net47 inh_ground_gnd3i inh_ground_gnd3i NE3I W=420.0n L=800n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM8 net035 net039 inh_ground_gnd3i inh_ground_gnd3i NE3I W=420.0n L=1u M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM7 net35 net039 net035 inh_ground_gnd3i NE3I W=420.0n L=1u M=1.0 AD=2.016e-13 
+ AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
MM3 net039 net47 net31 inh_ground_gnd3i NE3I W=420.0n L=800n M=1.0 
+ AD=2.016e-13 AS=2.016e-13 PD=1.8e-06 PS=1.8e-06 NRD=0.642857 NRS=0.642857
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    NA2I1JI3VX2
* View Name:    cmos_sch
************************************************************************

.SUBCKT NA2I1JI3VX2 AN B Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO AN:I B:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xnand2_1<0> B net4 Q inh_ground_gnd3i inh_power_vdd3i / nand2ji3v 
+ GT_PDL=350.00n GT_PDW=890.0n GT_PUL=300.00n GT_PUW=1.0u
Xnand2_1<1> B net4 Q inh_ground_gnd3i inh_power_vdd3i / nand2ji3v 
+ GT_PDL=350.00n GT_PDW=890.0n GT_PUL=300.00n GT_PUW=1.0u
Xinvr_1 AN net4 inh_ground_gnd3i inh_power_vdd3i / invrji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.41u
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    NA2JI3VX2
* View Name:    cmos_sch
************************************************************************

.SUBCKT NA2JI3VX2 A B Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xnand2_1<0> A B Q inh_ground_gnd3i inh_power_vdd3i / nand2ji3v GT_PDL=350.00n 
+ GT_PDW=890.0n GT_PUL=300.00n GT_PUW=1.00u
Xnand2_1<1> A B Q inh_ground_gnd3i inh_power_vdd3i / nand2ji3v GT_PDL=350.00n 
+ GT_PDW=890.0n GT_PUL=300.00n GT_PUW=1.00u
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    NO2JI3VX2
* View Name:    cmos_sch
************************************************************************

.SUBCKT NO2JI3VX2 A B Q inh_ground_gnd3i inh_power_vdd3i
*.PININFO A:I B:I Q:O inh_ground_gnd3i:B inh_power_vdd3i:B
Xnor2_1<0> A B Q inh_ground_gnd3i inh_power_vdd3i / nor2ji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.41u
Xnor2_1<1> A B Q inh_ground_gnd3i inh_power_vdd3i / nor2ji3v GT_PDL=350.00n 
+ GT_PDW=890.00n GT_PUL=300.00n GT_PUW=1.41u
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    DECAP5JI3V
* View Name:    cmos_sch
************************************************************************

.SUBCKT DECAP5JI3V inh_ground_gnd3i inh_power_vdd3i
*.PININFO inh_ground_gnd3i:B inh_power_vdd3i:B
MM0 net5 net4 inh_ground_gnd3i inh_ground_gnd3i NE3I W=830.0n L=1.48u M=1.0 
+ AD=3.984e-13 AS=3.984e-13 PD=2.62e-06 PS=2.62e-06 NRD=0.325301 NRS=0.325301
MM1 net4 net5 inh_power_vdd3i inh_power_vdd3i PE3I W=1.36u L=1.46u M=1.0 
+ AD=6.528e-13 AS=6.528e-13 PD=3.68e-06 PS=3.68e-06 NRD=0.198529 NRS=0.198529
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    DECAP7JI3V
* View Name:    cmos_sch
************************************************************************

.SUBCKT DECAP7JI3V inh_ground_gnd3i inh_power_vdd3i
*.PININFO inh_ground_gnd3i:B inh_power_vdd3i:B
MM7 net3 net4 inh_ground_gnd3i inh_ground_gnd3i NE3I W=880.0n L=350.0n M=1.0 
+ AD=4.224e-13 AS=4.224e-13 PD=2.72e-06 PS=2.72e-06 NRD=0.306818 NRS=0.306818
MM6 inh_ground_gnd3i net4 inh_ground_gnd3i inh_ground_gnd3i NE3I W=880.0n 
+ L=1.75u M=1.0 AD=4.224e-13 AS=4.224e-13 PD=2.72e-06 PS=2.72e-06 NRD=0.306818 
+ NRS=0.306818
MM5 net4 net3 inh_power_vdd3i inh_power_vdd3i PE3I W=1.315u L=300n M=1.0 
+ AD=6.312e-13 AS=6.312e-13 PD=3.59e-06 PS=3.59e-06 NRD=0.205323 NRS=0.205323
MM4 inh_power_vdd3i net3 inh_power_vdd3i inh_power_vdd3i PE3I W=1.315u L=1.71u 
+ M=1.0 AD=6.312e-13 AS=6.312e-13 PD=3.59e-06 PS=3.59e-06 NRD=0.205323 
+ NRS=0.205323
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    DECAP15JI3V
* View Name:    cmos_sch
************************************************************************

.SUBCKT DECAP15JI3V inh_ground_gnd3i inh_power_vdd3i
*.PININFO inh_ground_gnd3i:B inh_power_vdd3i:B
MM7 net3 net4 inh_ground_gnd3i inh_ground_gnd3i NE3I W=880.0n L=350.0n M=1.0 
+ AD=4.224e-13 AS=4.224e-13 PD=2.72e-06 PS=2.72e-06 NRD=0.306818 NRS=0.306818
MM6 inh_ground_gnd3i net4 inh_ground_gnd3i inh_ground_gnd3i NE3I W=2.64u 
+ L=1.71u M=1.0 AD=1.2672e-12 AS=1.2672e-12 PD=6.24e-06 PS=6.24e-06 
+ NRD=0.102273 NRS=0.102273
MM5 net4 net3 inh_power_vdd3i inh_power_vdd3i PE3I W=1.315u L=300n M=1.0 
+ AD=6.312e-13 AS=6.312e-13 PD=3.59e-06 PS=3.59e-06 NRD=0.205323 NRS=0.205323
MM4 inh_power_vdd3i net3 inh_power_vdd3i inh_power_vdd3i PE3I W=3.945u L=1.7u 
+ M=1.0 AD=1.8936e-12 AS=1.8936e-12 PD=8.85e-06 PS=8.85e-06 NRD=0.0684411 
+ NRS=0.0684411
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    DECAP25JI3V
* View Name:    cmos_sch
************************************************************************

.SUBCKT DECAP25JI3V inh_ground_gnd3i inh_power_vdd3i
*.PININFO inh_ground_gnd3i:B inh_power_vdd3i:B
MM7 net3 net4 inh_ground_gnd3i inh_ground_gnd3i NE3I W=880.0n L=350.0n M=1.0 
+ AD=4.224e-13 AS=4.224e-13 PD=2.72e-06 PS=2.72e-06 NRD=0.306818 NRS=0.306818
MM6 inh_ground_gnd3i net4 inh_ground_gnd3i inh_ground_gnd3i NE3I W=4.4u 
+ L=1.94u M=1.0 AD=2.112e-12 AS=2.112e-12 PD=9.76e-06 PS=9.76e-06 
+ NRD=0.0613636 NRS=0.0613636
MM5 net4 net3 inh_power_vdd3i inh_power_vdd3i PE3I W=1.315u L=300n M=1.0 
+ AD=6.312e-13 AS=6.312e-13 PD=3.59e-06 PS=3.59e-06 NRD=0.205323 NRS=0.205323
MM4 inh_power_vdd3i net3 inh_power_vdd3i inh_power_vdd3i PE3I W=6.575u L=1.93u 
+ M=1.0 AD=3.156e-12 AS=3.156e-12 PD=1.411e-05 PS=1.411e-05 NRD=0.0410646 
+ NRS=0.0410646
.ENDS

************************************************************************
* Library Name: D_CELLS_JI3V
* Cell Name:    DECAP10JI3V
* View Name:    cmos_sch
************************************************************************

.SUBCKT DECAP10JI3V inh_ground_gnd3i inh_power_vdd3i
*.PININFO inh_ground_gnd3i:B inh_power_vdd3i:B
MM7 net3 net4 inh_ground_gnd3i inh_ground_gnd3i NE3I W=880.0n L=350.0n M=1.0 
+ AD=4.224e-13 AS=4.224e-13 PD=2.72e-06 PS=2.72e-06 NRD=0.306818 NRS=0.306818
MM6 inh_ground_gnd3i net4 inh_ground_gnd3i inh_ground_gnd3i NE3I W=1.76u 
+ L=1.445u M=1.0 AD=8.448e-13 AS=8.448e-13 PD=4.48e-06 PS=4.48e-06 
+ NRD=0.153409 NRS=0.153409
MM5 net4 net3 inh_power_vdd3i inh_power_vdd3i PE3I W=1.315u L=300n M=1.0 
+ AD=6.312e-13 AS=6.312e-13 PD=3.59e-06 PS=3.59e-06 NRD=0.205323 NRS=0.205323
MM4 inh_power_vdd3i net3 inh_power_vdd3i inh_power_vdd3i PE3I W=2.63u L=1.425u 
+ M=1.0 AD=1.2624e-12 AS=1.2624e-12 PD=6.22e-06 PS=6.22e-06 NRD=0.102662 
+ NRS=0.102662
.ENDS

************************************************************************
* Library Name: ASKA_DIG2
* Cell Name:    aska_dig
* View Name:    schematic
************************************************************************

.SUBCKT aska_dig DAC<5> DAC<4> DAC<3> DAC<2> DAC<1> DAC<0> IC_addr<1> 
+ IC_addr<0> SPI_CS SPI_Clk SPI_MOSI clk down_switches<31> down_switches<30> 
+ down_switches<29> down_switches<28> down_switches<27> down_switches<26> 
+ down_switches<25> down_switches<24> down_switches<23> down_switches<22> 
+ down_switches<21> down_switches<20> down_switches<19> down_switches<18> 
+ down_switches<17> down_switches<16> down_switches<15> down_switches<14> 
+ down_switches<13> down_switches<12> down_switches<11> down_switches<10> 
+ down_switches<9> down_switches<8> down_switches<7> down_switches<6> 
+ down_switches<5> down_switches<4> down_switches<3> down_switches<2> 
+ down_switches<1> down_switches<0> enable porborn pulse_active reset_l 
+ up_switches<31> up_switches<30> up_switches<29> up_switches<28> 
+ up_switches<27> up_switches<26> up_switches<25> up_switches<24> 
+ up_switches<23> up_switches<22> up_switches<21> up_switches<20> 
+ up_switches<19> up_switches<18> up_switches<17> up_switches<16> 
+ up_switches<15> up_switches<14> up_switches<13> up_switches<12> 
+ up_switches<11> up_switches<10> up_switches<9> up_switches<8> up_switches<7> 
+ up_switches<6> up_switches<5> up_switches<4> up_switches<3> up_switches<2> 
+ up_switches<1> up_switches<0>
*.PININFO IC_addr<1>:I IC_addr<0>:I SPI_CS:I SPI_Clk:I SPI_MOSI:I clk:I 
*.PININFO porborn:I reset_l:I DAC<5>:O DAC<4>:O DAC<3>:O DAC<2>:O DAC<1>:O 
*.PININFO DAC<0>:O down_switches<31>:O down_switches<30>:O down_switches<29>:O 
*.PININFO down_switches<28>:O down_switches<27>:O down_switches<26>:O 
*.PININFO down_switches<25>:O down_switches<24>:O down_switches<23>:O 
*.PININFO down_switches<22>:O down_switches<21>:O down_switches<20>:O 
*.PININFO down_switches<19>:O down_switches<18>:O down_switches<17>:O 
*.PININFO down_switches<16>:O down_switches<15>:O down_switches<14>:O 
*.PININFO down_switches<13>:O down_switches<12>:O down_switches<11>:O 
*.PININFO down_switches<10>:O down_switches<9>:O down_switches<8>:O 
*.PININFO down_switches<7>:O down_switches<6>:O down_switches<5>:O 
*.PININFO down_switches<4>:O down_switches<3>:O down_switches<2>:O 
*.PININFO down_switches<1>:O down_switches<0>:O enable:O pulse_active:O 
*.PININFO up_switches<31>:O up_switches<30>:O up_switches<29>:O 
*.PININFO up_switches<28>:O up_switches<27>:O up_switches<26>:O 
*.PININFO up_switches<25>:O up_switches<24>:O up_switches<23>:O 
*.PININFO up_switches<22>:O up_switches<21>:O up_switches<20>:O 
*.PININFO up_switches<19>:O up_switches<18>:O up_switches<17>:O 
*.PININFO up_switches<16>:O up_switches<15>:O up_switches<14>:O 
*.PININFO up_switches<13>:O up_switches<12>:O up_switches<11>:O 
*.PININFO up_switches<10>:O up_switches<9>:O up_switches<8>:O up_switches<7>:O 
*.PININFO up_switches<6>:O up_switches<5>:O up_switches<4>:O up_switches<3>:O 
*.PININFO up_switches<2>:O up_switches<1>:O up_switches<0>:O
Xspi1_g992__7410 spi1_Rx_count<0> spi1_Rx_count<1> spi1_n_2018 gnd3i! vdd3i! / 
+ AND2JI3VX0
Xg17165 npg1_phase_down_state ele2<16> n_736 gnd3i! vdd3i! / AND2JI3VX0
Xg17163 npg1_phase_down_state ele2<31> n_734 gnd3i! vdd3i! / AND2JI3VX0
Xg17161 npg1_phase_down_state ele2<30> n_732 gnd3i! vdd3i! / AND2JI3VX0
Xg3 npg1_phase_down_state ele2<29> n_730 gnd3i! vdd3i! / AND2JI3VX0
Xg16922__2883 n_198 npg1_OFF_count<4> n_216 gnd3i! vdd3i! / AND2JI3VX0
Xg16915__1881 n_196 n_199 n_220 gnd3i! vdd3i! / AND2JI3VX0
Xg17167 n_180 n_108 n_739 gnd3i! vdd3i! / AND2JI3VX0
Xg17031__6783 FE_PHN233_npg1_OFF_count_3 conf1<13> n_112 gnd3i! vdd3i! / 
+ AND2JI3VX0
Xg17032__3680 n_38 conf0<7> n_111 gnd3i! vdd3i! / AND2JI3VX0
Xg16986__2883 n_97 n_101 n_163 gnd3i! vdd3i! / AND2JI3VX0
Xspi1_conf0_meta_reg[0] CTS_1 spi1_conf0_asyn<0> spi1_conf0_meta<0> 
+ FE_PHN263_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[1] CTS_1 spi1_conf0_asyn<1> spi1_conf0_meta<1> 
+ FE_PHN263_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[2] CTS_1 spi1_conf0_asyn<2> spi1_conf0_meta<2> 
+ FE_PHN263_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[3] CTS_1 spi1_conf0_asyn<3> spi1_conf0_meta<3> 
+ FE_PHN263_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[4] CTS_1 spi1_conf0_asyn<4> spi1_conf0_meta<4> 
+ FE_PHN263_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[5] CTS_1 spi1_conf0_asyn<5> spi1_conf0_meta<5> 
+ FE_PHN263_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[6] CTS_1 spi1_conf0_asyn<6> spi1_conf0_meta<6> 
+ FE_PHN263_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[7] CTS_1 spi1_conf0_asyn<7> spi1_conf0_meta<7> 
+ FE_PHN263_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[8] CTS_1 spi1_conf0_asyn<8> spi1_conf0_meta<8> 
+ FE_PHN263_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[9] CTS_1 spi1_conf0_asyn<9> spi1_conf0_meta<9> 
+ FE_PHN263_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[10] CTS_1 spi1_conf0_asyn<10> spi1_conf0_meta<10> 
+ FE_PHN263_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[11] CTS_1 spi1_conf0_asyn<11> spi1_conf0_meta<11> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[12] CTS_5 spi1_conf0_asyn<12> spi1_conf0_meta<12> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[13] CTS_5 spi1_conf0_asyn<13> spi1_conf0_meta<13> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[14] CTS_5 spi1_conf0_asyn<14> spi1_conf0_meta<14> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[15] CTS_5 spi1_conf0_asyn<15> spi1_conf0_meta<15> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[16] CTS_5 spi1_conf0_asyn<16> spi1_conf0_meta<16> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[17] CTS_2 spi1_conf0_asyn<17> spi1_conf0_meta<17> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[21] CTS_2 spi1_conf0_asyn<21> spi1_conf0_meta<21> 
+ FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[22] CTS_2 spi1_conf0_asyn<22> spi1_conf0_meta<22> 
+ FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[23] CTS_4 spi1_conf0_asyn<23> spi1_conf0_meta<23> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[24] CTS_4 spi1_conf0_asyn<24> spi1_conf0_meta<24> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[25] CTS_4 spi1_conf0_asyn<25> spi1_conf0_meta<25> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[26] CTS_4 spi1_conf0_asyn<26> spi1_conf0_meta<26> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[27] CTS_4 spi1_conf0_asyn<27> spi1_conf0_meta<27> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[28] CTS_4 spi1_conf0_asyn<28> spi1_conf0_meta<28> 
+ FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[29] CTS_4 spi1_conf0_asyn<29> spi1_conf0_meta<29> 
+ FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[30] CTS_4 spi1_conf0_asyn<30> spi1_conf0_meta<30> 
+ FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[31] CTS_4 spi1_conf0_asyn<31> spi1_conf0_meta<31> 
+ FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[0] CTS_1 spi1_conf1_asyn<0> spi1_conf1_meta<0> 
+ FE_PHN263_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[2] CTS_1 spi1_conf1_asyn<2> spi1_conf1_meta<2> 
+ FE_PHN263_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[4] CTS_1 spi1_conf1_asyn<4> spi1_conf1_meta<4> 
+ FE_PHN263_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[5] CTS_1 spi1_conf1_asyn<5> spi1_conf1_meta<5> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[6] CTS_1 spi1_conf1_asyn<6> spi1_conf1_meta<6> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[7] CTS_1 spi1_conf1_asyn<7> spi1_conf1_meta<7> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[8] CTS_1 spi1_conf1_asyn<8> spi1_conf1_meta<8> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[9] CTS_1 spi1_conf1_asyn<9> spi1_conf1_meta<9> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[14] CTS_5 spi1_conf1_asyn<14> spi1_conf1_meta<14> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[15] CTS_2 spi1_conf1_asyn<15> spi1_conf1_meta<15> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[16] CTS_2 spi1_conf1_asyn<16> spi1_conf1_meta<16> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[17] CTS_5 spi1_conf1_asyn<17> spi1_conf1_meta<17> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[18] CTS_2 spi1_conf1_asyn<18> spi1_conf1_meta<18> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[19] CTS_2 spi1_conf1_asyn<19> spi1_conf1_meta<19> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[20] CTS_2 spi1_conf1_asyn<20> spi1_conf1_meta<20> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[21] CTS_4 spi1_conf1_asyn<21> spi1_conf1_meta<21> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[22] CTS_4 spi1_conf1_asyn<22> spi1_conf1_meta<22> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[23] CTS_4 spi1_conf1_asyn<23> spi1_conf1_meta<23> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[0] CTS_5 spi1_ele1_asyn<0> spi1_ele1_meta<0> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[1] CTS_1 spi1_ele1_asyn<1> spi1_ele1_meta<1> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[2] CTS_1 spi1_ele1_asyn<2> spi1_ele1_meta<2> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[3] CTS_1 spi1_ele1_asyn<3> spi1_ele1_meta<3> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[4] CTS_1 spi1_ele1_asyn<4> spi1_ele1_meta<4> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[5] CTS_1 spi1_ele1_asyn<5> spi1_ele1_meta<5> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[6] CTS_1 spi1_ele1_asyn<6> spi1_ele1_meta<6> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[7] CTS_1 spi1_ele1_asyn<7> spi1_ele1_meta<7> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[8] CTS_1 spi1_ele1_asyn<8> spi1_ele1_meta<8> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[9] CTS_5 spi1_ele1_asyn<9> spi1_ele1_meta<9> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[10] CTS_5 spi1_ele1_asyn<10> spi1_ele1_meta<10> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[11] CTS_5 spi1_ele1_asyn<11> spi1_ele1_meta<11> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[12] CTS_5 spi1_ele1_asyn<12> spi1_ele1_meta<12> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[15] CTS_5 spi1_ele1_asyn<15> spi1_ele1_meta<15> 
+ FE_OFN35_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[16] CTS_5 spi1_ele1_asyn<16> spi1_ele1_meta<16> 
+ FE_OFN35_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[17] CTS_5 spi1_ele1_asyn<17> spi1_ele1_meta<17> 
+ FE_OFN35_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[18] CTS_5 spi1_ele1_asyn<18> spi1_ele1_meta<18> 
+ FE_OFN35_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[19] CTS_5 spi1_ele1_asyn<19> spi1_ele1_meta<19> 
+ FE_OFN35_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[20] CTS_5 spi1_ele1_asyn<20> spi1_ele1_meta<20> 
+ FE_OFN35_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[21] CTS_5 spi1_ele1_asyn<21> spi1_ele1_meta<21> 
+ FE_OFN35_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[22] CTS_5 spi1_ele1_asyn<22> spi1_ele1_meta<22> 
+ FE_OFN35_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[23] CTS_4 spi1_ele1_asyn<23> spi1_ele1_meta<23> 
+ FE_OFN35_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[24] CTS_4 spi1_ele1_asyn<24> spi1_ele1_meta<24> 
+ FE_OFN35_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[25] CTS_4 spi1_ele1_asyn<25> spi1_ele1_meta<25> 
+ FE_OFN35_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[26] CTS_4 spi1_ele1_asyn<26> spi1_ele1_meta<26> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[27] CTS_4 spi1_ele1_asyn<27> spi1_ele1_meta<27> 
+ FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[28] CTS_4 spi1_ele1_asyn<28> spi1_ele1_meta<28> 
+ FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[29] CTS_4 spi1_ele1_asyn<29> spi1_ele1_meta<29> 
+ FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[30] CTS_4 spi1_ele1_asyn<30> spi1_ele1_meta<30> 
+ FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[31] CTS_4 spi1_ele1_asyn<31> spi1_ele1_meta<31> 
+ FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[0] CTS_5 spi1_ele2_asyn<0> spi1_ele2_meta<0> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[1] CTS_1 spi1_ele2_asyn<1> spi1_ele2_meta<1> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[2] CTS_1 spi1_ele2_asyn<2> spi1_ele2_meta<2> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[3] CTS_1 spi1_ele2_asyn<3> spi1_ele2_meta<3> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[4] CTS_1 spi1_ele2_asyn<4> spi1_ele2_meta<4> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[5] CTS_1 spi1_ele2_asyn<5> spi1_ele2_meta<5> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[6] CTS_1 spi1_ele2_asyn<6> spi1_ele2_meta<6> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[7] CTS_1 spi1_ele2_asyn<7> spi1_ele2_meta<7> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[8] CTS_1 spi1_ele2_asyn<8> spi1_ele2_meta<8> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[9] CTS_5 spi1_ele2_asyn<9> spi1_ele2_meta<9> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[10] CTS_5 spi1_ele2_asyn<10> spi1_ele2_meta<10> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[11] CTS_5 spi1_ele2_asyn<11> spi1_ele2_meta<11> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[12] CTS_5 spi1_ele2_asyn<12> spi1_ele2_meta<12> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[14] CTS_5 spi1_ele2_asyn<14> spi1_ele2_meta<14> 
+ FE_OFN35_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[15] CTS_5 spi1_ele2_asyn<15> spi1_ele2_meta<15> 
+ FE_OFN35_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[16] CTS_5 spi1_ele2_asyn<16> spi1_ele2_meta<16> 
+ FE_OFN35_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[17] CTS_5 spi1_ele2_asyn<17> spi1_ele2_meta<17> 
+ FE_OFN35_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[18] CTS_5 spi1_ele2_asyn<18> spi1_ele2_meta<18> 
+ FE_OFN35_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[19] CTS_5 spi1_ele2_asyn<19> spi1_ele2_meta<19> 
+ FE_OFN35_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[20] CTS_5 spi1_ele2_asyn<20> spi1_ele2_meta<20> 
+ FE_OFN35_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[21] CTS_5 spi1_ele2_asyn<21> spi1_ele2_meta<21> 
+ FE_OFN35_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[22] CTS_5 spi1_ele2_asyn<22> spi1_ele2_meta<22> 
+ FE_OFN35_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[23] CTS_4 spi1_ele2_asyn<23> spi1_ele2_meta<23> 
+ FE_OFN35_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[24] CTS_4 spi1_ele2_asyn<24> spi1_ele2_meta<24> 
+ FE_OFN35_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[25] CTS_4 spi1_ele2_asyn<25> spi1_ele2_meta<25> 
+ FE_OFN35_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[26] CTS_4 spi1_ele2_asyn<26> spi1_ele2_meta<26> 
+ FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[27] CTS_4 spi1_ele2_asyn<27> spi1_ele2_meta<27> 
+ FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[28] CTS_4 spi1_ele2_asyn<28> spi1_ele2_meta<28> 
+ FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[29] CTS_4 spi1_ele2_asyn<29> spi1_ele2_meta<29> 
+ FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[30] CTS_4 spi1_ele2_asyn<30> spi1_ele2_meta<30> 
+ FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_UP_accumulator_reg[0] CTS_1 n_454 npg1_UP_accumulator<0> FE_PHN440_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_UP_accumulator_reg[1] CTS_1 n_453 npg1_UP_accumulator<1> FE_PHN441_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_UP_accumulator_reg[2] CTS_1 n_452 npg1_UP_accumulator<2> FE_PHN263_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_UP_accumulator_reg[3] CTS_1 n_451 npg1_UP_accumulator<3> FE_PHN433_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_UP_accumulator_reg[4] CTS_1 n_450 npg1_UP_accumulator<4> FE_PHN434_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_UP_accumulator_reg[5] CTS_2 n_482 npg1_UP_accumulator<5> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_UP_accumulator_reg[6] CTS_1 n_490 npg1_UP_accumulator<6> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_UP_accumulator_reg[7] CTS_2 n_495 npg1_UP_accumulator<7> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_UP_accumulator_reg[8] CTS_2 n_503 npg1_UP_accumulator<8> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_UP_accumulator_reg[9] CTS_2 n_506 npg1_UP_accumulator<9> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_Rx_count_reg[5] CTS_8 FE_PHN410_spi1_n_1763 spi1_Rx_count<5> 
+ FE_OFN30_SPI_CS gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_Rx_count_reg[4] CTS_8 spi1_n_1924 spi1_Rx_count<4> FE_OFN30_SPI_CS 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_Rx_count_reg[3] CTS_8 spi1_n_1962 spi1_Rx_count<3> FE_OFN30_SPI_CS 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_on_off_ctrl_reg[2] CTS_2 n_302 npg1_on_off_ctrl<2> FE_PHN442_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_on_off_ctrl_reg[1] CTS_2 n_306 npg1_on_off_ctrl<1> FE_PHN436_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[1] CTS_1 FE_PHN348_spi1_conf1_meta_1 conf1<1> FE_PHN439_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[3] CTS_1 FE_PHN293_spi1_conf1_meta_3 conf1<3> FE_PHN435_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[6] CTS_1 FE_PHN303_spi1_conf1_meta_6 conf1<6> FE_PHN432_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_Rx_count_reg[1] CTS_8 spi1_n_2008 spi1_Rx_count<1> FE_OFN30_SPI_CS 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[31] CTS_4 FE_PHN296_spi1_ele2_meta_31 ele2<31> FE_PHN271_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[30] CTS_4 FE_PHN338_spi1_ele2_meta_30 ele2<30> FE_PHN271_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[29] CTS_4 FE_PHN276_spi1_ele2_meta_29 ele2<29> FE_PHN271_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[28] CTS_4 FE_PHN333_spi1_ele2_meta_28 ele2<28> FE_PHN271_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[27] CTS_4 FE_PHN340_spi1_ele2_meta_27 ele2<27> FE_PHN431_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[13] CTS_2 spi1_conf1_asyn<13> spi1_conf1_meta<13> 
+ FE_PHN444_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[19] CTS_2 spi1_conf0_asyn<19> spi1_conf0_meta<19> 
+ FE_PHN443_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[1] CTS_1 spi1_conf1_asyn<1> spi1_conf1_meta<1> 
+ FE_PHN438_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[3] CTS_1 spi1_conf1_asyn<3> spi1_conf1_meta<3> 
+ FE_PHN437_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[10] CTS_2 spi1_conf1_asyn<10> spi1_conf1_meta<10> 
+ FE_PHN446_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[11] CTS_2 spi1_conf1_asyn<11> spi1_conf1_meta<11> 
+ FE_PHN446_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_meta_reg[12] CTS_2 spi1_conf1_asyn<12> spi1_conf1_meta<12> 
+ FE_PHN446_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[18] CTS_2 spi1_conf0_asyn<18> spi1_conf0_meta<18> 
+ FE_PHN446_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_meta_reg[20] CTS_2 spi1_conf0_asyn<20> spi1_conf0_meta<20> 
+ FE_PHN446_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_DOWN_accumulator_reg[0] CTS_2 n_383 npg1_DOWN_accumulator<0> 
+ FE_PHN447_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_DOWN_accumulator_reg[1] CTS_2 n_382 npg1_DOWN_accumulator<1> 
+ FE_PHN447_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_DOWN_accumulator_reg[2] CTS_2 n_381 npg1_DOWN_accumulator<2> 
+ FE_PHN445_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_DOWN_accumulator_reg[3] CTS_2 n_402 npg1_DOWN_accumulator<3> 
+ FE_PHN445_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_DOWN_accumulator_reg[4] CTS_2 n_434 npg1_DOWN_accumulator<4> 
+ FE_PHN445_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_DOWN_accumulator_reg[5] CTS_2 n_483 npg1_DOWN_accumulator<5> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_DOWN_accumulator_reg[6] CTS_2 n_489 npg1_DOWN_accumulator<6> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_DOWN_accumulator_reg[7] CTS_2 n_496 npg1_DOWN_accumulator<7> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_DOWN_accumulator_reg[8] CTS_2 n_504 npg1_DOWN_accumulator<8> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_DOWN_accumulator_reg[9] CTS_2 n_505 npg1_DOWN_accumulator<9> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[20] CTS_2 FE_PHN366_spi1_conf0_meta_20 conf0<20> 
+ FE_PHN446_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[19] CTS_2 FE_PHN346_spi1_conf0_meta_19 conf0<19> 
+ FE_PHN446_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[5] CTS_2 FE_PHN396_spi1_conf1_meta_5 conf1<5> FE_PHN445_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[8] CTS_5 FE_PHN395_spi1_ele2_meta_8 ele2<8> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[9] CTS_2 FE_PHN394_spi1_conf1_meta_9 conf1<9> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[6] CTS_1 FE_PHN393_spi1_ele2_meta_6 ele2<6> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[8] CTS_5 FE_PHN392_spi1_ele1_meta_8 ele1<8> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[19] CTS_5 FE_PHN391_spi1_ele1_meta_19 ele1<19> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[21] CTS_2 FE_PHN390_spi1_conf0_meta_21 conf0<21> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[7] CTS_2 FE_PHN389_spi1_conf1_meta_7 conf1<7> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[26] CTS_4 FE_PHN388_spi1_ele2_meta_26 ele2<26> FE_PHN431_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[4] CTS_1 FE_PHN387_spi1_conf1_meta_4 conf1<4> FE_PHN263_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[0] CTS_1 FE_PHN386_spi1_conf0_meta_0 conf0<0> FE_PHN263_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[14] CTS_5 FE_PHN385_spi1_ele2_meta_14 ele2<14> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[16] CTS_2 FE_PHN384_spi1_conf1_meta_16 conf1<16> FE_OFN33_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[22] CTS_5 FE_PHN383_spi1_ele2_meta_22 ele2<22> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[2] CTS_1 FE_PHN382_spi1_ele1_meta_2 ele1<2> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[24] CTS_4 FE_PHN381_spi1_ele1_meta_24 ele1<24> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[10] CTS_5 FE_PHN380_spi1_ele2_meta_10 ele2<10> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[30] CTS_4 FE_PHN379_spi1_conf0_meta_30 conf0<30> 
+ FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[17] CTS_2 FE_PHN378_spi1_conf1_meta_17 conf1<17> FE_OFN33_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[18] CTS_2 FE_PHN377_spi1_conf0_meta_18 conf0<18> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[2] CTS_1 FE_PHN376_spi1_conf1_meta_2 conf1<2> FE_PHN263_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[31] CTS_4 FE_PHN375_spi1_ele1_meta_31 ele1<31> FE_PHN271_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[10] CTS_2 FE_PHN374_spi1_conf1_meta_10 conf1<10> FE_OFN33_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[27] CTS_4 FE_PHN373_spi1_conf0_meta_27 conf0<27> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[12] CTS_2 FE_PHN372_spi1_conf1_meta_12 conf1<12> FE_OFN33_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[29] CTS_4 FE_PHN371_spi1_ele1_meta_29 ele1<29> FE_PHN271_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[16] CTS_5 FE_PHN370_spi1_ele1_meta_16 ele1<16> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[5] CTS_1 FE_PHN369_spi1_conf0_meta_5 conf0<5> FE_PHN263_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[16] CTS_5 FE_PHN368_spi1_ele2_meta_16 ele2<16> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[8] CTS_1 FE_PHN367_spi1_conf0_meta_8 conf0<8> FE_PHN263_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[13] CTS_5 FE_PHN365_spi1_conf0_meta_13 conf0<13> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[24] CTS_4 FE_PHN364_spi1_conf0_meta_24 conf0<24> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[22] CTS_5 FE_PHN363_spi1_ele1_meta_22 ele1<22> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[28] CTS_4 FE_PHN362_spi1_ele1_meta_28 ele1<28> FE_PHN271_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[11] CTS_2 FE_PHN361_spi1_conf1_meta_11 conf1<11> FE_OFN33_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[14] CTS_5 FE_PHN360_spi1_conf0_meta_14 conf0<14> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[23] CTS_4 FE_PHN359_spi1_ele1_meta_23 ele1<23> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[7] CTS_1 FE_PHN358_spi1_ele2_meta_7 ele2<7> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[9] CTS_1 FE_PHN357_spi1_conf0_meta_9 conf0<9> FE_PHN263_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[21] CTS_4 FE_PHN356_spi1_conf1_meta_21 conf1<21> 
+ FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[23] CTS_4 FE_PHN355_spi1_conf1_meta_23 conf1<23> 
+ FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[17] CTS_5 FE_PHN354_spi1_ele1_meta_17 ele1<17> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[7] CTS_1 FE_PHN353_spi1_conf0_meta_7 conf0<7> FE_PHN263_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[22] CTS_4 FE_PHN352_spi1_conf1_meta_22 conf1<22> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[13] CTS_2 FE_PHN351_spi1_conf1_meta_13 conf1<13> FE_OFN33_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[6] CTS_1 FE_PHN350_spi1_ele1_meta_6 ele1<6> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[0] CTS_5 FE_PHN349_spi1_ele1_meta_0 ele1<0> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[26] CTS_4 FE_PHN347_spi1_conf0_meta_26 conf0<26> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[22] CTS_2 FE_PHN298_spi1_conf0_meta_22 conf0<22> FE_OFN33_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_phase_up_state_reg CTS_4 n_281 npg1_phase_up_state FE_PHN271_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[28] CTS_4 FE_PHN345_spi1_conf0_meta_28 conf0<28> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[26] CTS_4 FE_PHN344_spi1_ele1_meta_26 ele1<26> FE_PHN431_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[3] CTS_1 FE_PHN343_spi1_ele2_meta_3 ele2<3> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[25] CTS_4 FE_PHN342_spi1_conf0_meta_25 conf0<25> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[15] CTS_5 FE_PHN341_spi1_ele2_meta_15 ele2<15> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[7] CTS_1 FE_PHN337_spi1_ele1_meta_7 ele1<7> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[24] CTS_4 FE_PHN336_spi1_ele2_meta_24 ele2<24> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[30] CTS_4 FE_PHN335_spi1_ele1_meta_30 ele1<30> FE_PHN271_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[6] CTS_1 FE_PHN334_spi1_conf0_meta_6 conf0<6> FE_PHN263_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[5] CTS_1 FE_PHN332_spi1_ele1_meta_5 ele1<5> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[12] CTS_5 FE_PHN331_spi1_ele2_meta_12 ele2<12> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[1] CTS_1 FE_PHN330_spi1_ele1_meta_1 ele1<1> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[20] CTS_5 FE_PHN328_spi1_ele1_meta_20 ele1<20> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[25] CTS_4 FE_PHN327_spi1_ele1_meta_25 ele1<25> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[4] CTS_1 FE_PHN326_spi1_ele1_meta_4 ele1<4> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[11] CTS_5 FE_PHN325_spi1_ele2_meta_11 ele2<11> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[2] CTS_1 FE_PHN324_spi1_ele2_meta_2 ele2<2> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[13] CTS_5 FE_PHN323_spi1_ele1_meta_13 ele1<13> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[3] CTS_1 FE_PHN322_spi1_ele1_meta_3 ele1<3> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[18] CTS_5 FE_PHN321_spi1_ele1_meta_18 ele1<18> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[5] CTS_1 FE_PHN320_spi1_ele2_meta_5 ele2<5> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[23] CTS_4 FE_PHN319_spi1_ele2_meta_23 ele2<23> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[29] CTS_4 FE_PHN318_spi1_conf0_meta_29 conf0<29> 
+ FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[12] CTS_5 FE_PHN317_spi1_conf0_meta_12 conf0<12> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[21] CTS_5 FE_PHN316_spi1_ele1_meta_21 ele1<21> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[20] CTS_5 FE_PHN315_spi1_ele2_meta_20 ele2<20> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[25] CTS_4 FE_PHN313_spi1_ele2_meta_25 ele2<25> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[13] CTS_5 FE_PHN312_spi1_ele2_meta_13 ele2<13> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[21] CTS_5 FE_PHN311_spi1_ele2_meta_21 ele2<21> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[10] CTS_1 FE_PHN310_spi1_conf0_meta_10 conf0<10> 
+ FE_PHN263_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[27] CTS_4 FE_PHN309_spi1_ele1_meta_27 ele1<27> FE_PHN431_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[9] CTS_5 FE_PHN308_spi1_ele1_meta_9 ele1<9> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[17] CTS_2 FE_PHN307_spi1_conf0_meta_17 conf0<17> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[19] CTS_5 FE_PHN306_spi1_ele2_meta_19 ele2<19> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[1] CTS_1 FE_PHN305_spi1_conf0_meta_1 conf0<1> FE_PHN263_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[16] CTS_5 FE_PHN304_spi1_conf0_meta_16 conf0<16> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[23] CTS_4 FE_PHN302_spi1_conf0_meta_23 conf0<23> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[15] CTS_5 FE_PHN301_spi1_ele1_meta_15 ele1<15> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[9] CTS_5 FE_PHN300_spi1_ele2_meta_9 ele2<9> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[1] CTS_1 FE_PHN299_spi1_ele2_meta_1 ele2<1> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[10] CTS_5 FE_PHN297_spi1_ele1_meta_10 ele1<10> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[18] CTS_5 FE_PHN295_spi1_ele2_meta_18 ele2<18> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[0] CTS_5 FE_PHN290_spi1_ele2_meta_0 ele2<0> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[4] CTS_1 FE_PHN289_spi1_ele2_meta_4 ele2<4> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[31] CTS_4 FE_PHN288_spi1_conf0_meta_31 conf0<31> 
+ FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[15] CTS_5 FE_PHN286_spi1_conf0_meta_15 conf0<15> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[14] CTS_5 FE_PHN285_spi1_ele1_meta_14 ele1<14> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[3] CTS_1 FE_PHN284_spi1_conf0_meta_3 conf0<3> FE_PHN263_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[2] CTS_1 FE_PHN283_spi1_conf0_meta_2 conf0<2> FE_PHN263_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[4] CTS_1 FE_PHN281_spi1_conf0_meta_4 conf0<4> FE_PHN263_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf0_reg[11] CTS_1 FE_PHN280_spi1_conf0_meta_11 conf0<11> 
+ FE_PHN263_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_reg[17] CTS_5 FE_PHN279_spi1_ele2_meta_17 ele2<17> FE_OFN35_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[12] CTS_5 FE_PHN278_spi1_ele1_meta_12 ele1<12> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_reg[11] CTS_5 FE_PHN277_spi1_ele1_meta_11 ele1<11> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_phase_down_state_reg CTS_4 n_738 npg1_phase_down_state FE_PHN271_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_DOWN_count_reg[5] CTS_2 n_410 npg1_DOWN_count<5> FE_OFN33_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_OFF_count_reg[0] CTS_2 n_441 npg1_OFF_count<0> FE_OFN33_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_OFF_count_reg[5] CTS_2 n_436 npg1_OFF_count<5> FE_OFN33_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_OFF_count_reg[6] CTS_2 n_439 npg1_OFF_count<6> FE_OFN33_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_OFF_count_reg[4] CTS_2 n_469 npg1_OFF_count<4> FE_OFN33_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_on_off_ctrl_reg[0] CTS_2 n_336 npg1_on_off_ctrl<0> FE_OFN33_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_DAC_cont_reg[0] CTS_5 n_349 npg1_DAC_cont<0> FE_OFN443_FE_PHN271_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[0] CTS_1 FE_PHN292_spi1_conf1_meta_0 conf1<0> FE_PHN263_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[8] CTS_1 FE_PHN329_spi1_conf1_meta_8 conf1<8> 
+ FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_OFF_count_reg[8] CTS_2 n_475 npg1_OFF_count<8> FE_OFN33_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_OFF_count_reg[7] CTS_2 n_438 npg1_OFF_count<7> FE_OFN33_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_OFF_count_reg[1] CTS_2 n_477 npg1_OFF_count<1> FE_OFN33_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_OFF_count_reg[2] CTS_2 n_468 npg1_OFF_count<2> FE_OFN33_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_OFF_count_reg[3] CTS_2 n_476 npg1_OFF_count<3> FE_OFN33_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[18] CTS_2 FE_PHN339_spi1_conf1_meta_18 conf1<18> FE_OFN33_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[19] CTS_2 FE_PHN294_spi1_conf1_meta_19 conf1<19> FE_OFN33_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[15] CTS_2 FE_PHN314_spi1_conf1_meta_15 conf1<15> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_freq_count_reg[8] CTS_1 n_408 npg1_freq_count<8> FE_PHN263_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_freq_count_reg[2] CTS_1 n_379 npg1_freq_count<2> FE_PHN263_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_freq_count_reg[10] CTS_1 n_429 npg1_freq_count<10> FE_PHN263_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_freq_count_reg[11] CTS_1 FE_PHN409_n_442 npg1_freq_count<11> 
+ FE_PHN263_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_freq_count_reg[4] CTS_1 n_380 npg1_freq_count<4> FE_PHN263_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_ON_count_reg[6] CTS_4 n_474 npg1_ON_count<6> FE_PHN271_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_ON_count_reg[5] CTS_4 n_435 npg1_ON_count<5> FE_PHN271_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_ON_count_reg[3] CTS_4 n_478 npg1_ON_count<3> FE_PHN431_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_ON_count_reg[4] CTS_4 n_470 npg1_ON_count<4> FE_PHN431_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_ON_count_reg[1] CTS_4 n_437 npg1_ON_count<1> FE_PHN431_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_ON_count_reg[2] CTS_4 n_440 npg1_ON_count<2> FE_PHN431_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_pulse_start_reg CTS_4 FE_PHN291_npg1_pulse_aux npg1_pulse_start 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_pulse_aux_reg CTS_4 n_276 npg1_pulse_aux FE_PHN431_n_32 gnd3i! vdd3i! / 
+ DFRRQJI3VX1
Xnpg1_freq_count_reg[7] CTS_1 n_398 npg1_freq_count<7> FE_PHN263_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_freq_count_reg[1] CTS_1 n_392 npg1_freq_count<1> FE_PHN263_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_freq_count_reg[5] CTS_1 n_354 npg1_freq_count<5> FE_PHN263_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_freq_count_reg[6] CTS_1 n_370 npg1_freq_count<6> FE_PHN263_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_phase_up_count_reg[0] CTS_4 n_299 npg1_phase_up_count<0> FE_PHN271_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_freq_count_reg[0] CTS_1 n_352 npg1_freq_count<0> FE_PHN263_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_freq_count_reg[3] CTS_1 n_389 npg1_freq_count<3> FE_PHN263_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_freq_count_reg[9] CTS_1 n_409 npg1_freq_count<9> FE_PHN263_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_UP_count_reg[4] CTS_2 n_484 npg1_UP_count<4> FE_PHN446_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_UP_count_reg[5] CTS_2 n_481 npg1_UP_count<5> FE_PHN446_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[20] CTS_2 FE_PHN287_spi1_conf1_meta_20 FE_OFN52_enable 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_conf1_reg[14] CTS_2 FE_PHN282_spi1_conf1_meta_14 conf1<14> 
+ FE_PHN431_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_DOWN_count_reg[4] CTS_2 n_412 npg1_DOWN_count<4> FE_PHN447_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_DOWN_count_reg[1] CTS_2 n_378 npg1_DOWN_count<1> FE_PHN447_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_DOWN_count_reg[2] CTS_2 n_385 npg1_DOWN_count<2> FE_PHN447_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_DOWN_count_reg[3] CTS_2 n_384 npg1_DOWN_count<3> FE_PHN447_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_UP_count_reg[1] CTS_2 n_449 npg1_UP_count<1> FE_PHN447_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_UP_count_reg[3] CTS_2 n_456 npg1_UP_count<3> FE_PHN447_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_UP_count_reg[2] CTS_2 n_448 npg1_UP_count<2> FE_PHN447_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX1
Xnpg1_DAC_cont_reg[5] CTS_5 n_471 npg1_DAC_cont<5> FE_PHN272_FE_OFN33_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_DAC_cont_reg[1] CTS_5 n_350 npg1_DAC_cont<1> FE_PHN272_FE_OFN33_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_DAC_cont_reg[2] CTS_5 FE_PHN411_n_391 npg1_DAC_cont<2> 
+ FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_DAC_cont_reg[4] CTS_5 n_455 npg1_DAC_cont<4> FE_PHN272_FE_OFN33_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_DAC_cont_reg[3] CTS_5 n_411 npg1_DAC_cont<3> FE_PHN272_FE_OFN33_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX1
Xnpg1_phase_down_count_reg[1] CTS_4 n_318 npg1_phase_down_count<1> 
+ FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[31] CTS_4 spi1_ele2_asyn<31> spi1_ele2_meta<31> 
+ FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele2_meta_reg[13] CTS_5 spi1_ele2_asyn<13> spi1_ele2_meta<13> 
+ FE_PHN446_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[13] CTS_5 spi1_ele1_asyn<13> spi1_ele1_meta<13> 
+ FE_PHN446_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_ele1_meta_reg[14] CTS_5 spi1_ele1_asyn<14> spi1_ele1_meta<14> 
+ FE_PHN446_n_32 gnd3i! vdd3i! / DFRRQJI3VX1
Xspi1_g986__9315 spi1_n_2017 spi1_n_2018 spi1_n_2008 gnd3i! vdd3i! / NO2JI3VX0
Xspi1_g991__1666 FE_PHN406_spi1_Rx_count_1 spi1_Rx_count<0> spi1_n_2017 gnd3i! 
+ vdd3i! / NO2JI3VX0
Xg11751__5115 FE_OFN15_up_switches_16 FE_OFN14_up_switches_17 n_637 gnd3i! 
+ vdd3i! / NO2JI3VX0
Xg11752__7482 FE_OFN2_up_switches_30 FE_OFN1_up_switches_31 n_636 gnd3i! 
+ vdd3i! / NO2JI3VX0
Xg11753__4733 FE_OFN4_up_switches_28 FE_OFN3_up_switches_29 n_635 gnd3i! 
+ vdd3i! / NO2JI3VX0
Xg11754__6161 FE_OFN13_up_switches_18 FE_OFN12_up_switches_19 n_634 gnd3i! 
+ vdd3i! / NO2JI3VX0
Xg16952__9945 FE_PHN233_npg1_OFF_count_3 n_159 n_198 gnd3i! vdd3i! / NO2JI3VX0
Xg16918__4733 n_169 n_182 n_217 gnd3i! vdd3i! / NO2JI3VX0
Xg17050__9315 conf0<12> n_25 n_96 gnd3i! vdd3i! / NO2JI3VX0
Xg16670__2398 n_403 n_432 n_446 gnd3i! vdd3i! / NO2JI3VX0
Xg16692__1881 npg1_OFF_count<0> n_414 n_432 gnd3i! vdd3i! / NO2JI3VX0
Xg16993__2398 npg1_on_off_ctrl<1> n_114 n_158 gnd3i! vdd3i! / NO2JI3VX0
Xg17080__7482 n_49 n_44 n_69 gnd3i! vdd3i! / NO2JI3VX0
Xg17081__4733 npg1_on_off_ctrl<2> npg1_on_off_ctrl<0> n_68 gnd3i! vdd3i! / 
+ NO2JI3VX0
Xg17056__9945 npg1_freq_count<2> n_35 n_60 gnd3i! vdd3i! / NO2JI3VX0
Xg16953__2883 n_42 n_135 n_197 gnd3i! vdd3i! / NO2JI3VX0
Xg16835__8428 n_16 n_289 n_304 gnd3i! vdd3i! / NO2JI3VX0
Xg16773__6131 n_38 n_313 n_362 gnd3i! vdd3i! / NO2JI3VX0
Xg16898__2398 npg1_pulse_start n_739 n_244 gnd3i! vdd3i! / NO2JI3VX0
Xg17069__6783 conf1<22> n_51 n_83 gnd3i! vdd3i! / NO2JI3VX0
Xg16803__2802 npg1_freq_count<0> n_320 n_340 gnd3i! vdd3i! / NO2JI3VX0
Xg16772__7098 n_11 n_340 n_364 gnd3i! vdd3i! / NO2JI3VX0
Xg17058__2346 npg1_UP_count<1> npg1_UP_count<0> n_58 gnd3i! vdd3i! / NO2JI3VX0
Xg16833__6260 n_124 n_269 n_305 gnd3i! vdd3i! / NO2JI3VX0
Xg17040__8246 conf0<1> n_35 n_106 gnd3i! vdd3i! / NO2JI3VX0
Xg17087__2346 n_55 npg1_UP_count<4> n_63 gnd3i! vdd3i! / NO2JI3VX0
Xg17088__1666 conf0<19> n_21 n_62 gnd3i! vdd3i! / NO2JI3VX0
Xg17047__4733 conf0<4> n_17 n_99 gnd3i! vdd3i! / NO2JI3VX0
Xg17025__2398 conf1<11> n_49 n_118 gnd3i! vdd3i! / NO2JI3VX0
Xg17079__5115 conf0<28> n_16 n_70 gnd3i! vdd3i! / NO2JI3VX0
Xg17046__7482 conf0<29> n_41 n_100 gnd3i! vdd3i! / NO2JI3VX0
Xg16882__6131 npg1_phase_down_count<1> n_243 n_254 gnd3i! vdd3i! / NO2JI3VX0
Xg17039__5122 conf1<14> n_50 n_107 gnd3i! vdd3i! / NO2JI3VX0
Xg17026__5107 conf1<13> FE_PHN233_npg1_OFF_count_3 n_117 gnd3i! vdd3i! / 
+ NO2JI3VX0
Xg17068__5526 conf1<15> n_46 n_84 gnd3i! vdd3i! / NO2JI3VX0
Xg16900__6260 npg1_phase_pause_ready n_214 n_243 gnd3i! vdd3i! / NO2JI3VX0
Xg17041__7098 conf0<8> n_15 n_104 gnd3i! vdd3i! / NO2JI3VX0
Xg16980__7482 n_99 n_74 n_151 gnd3i! vdd3i! / NO2JI3VX0
Xg17076__7098 conf0<5> n_52 n_74 gnd3i! vdd3i! / NO2JI3VX0
Xg17082__6161 conf0<9> n_36 n_67 gnd3i! vdd3i! / NO2JI3VX0
Xg17071__1617 conf0<10> n_54 n_81 gnd3i! vdd3i! / NO2JI3VX0
Xspi1_g939__1881 spi1_n_1998 spi1_Rx_data_temp<32> spi1_n_1994 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11881__2398 FE_PHN419_porborn reset_l npg1_n_374 gnd3i! vdd3i! / NA2JI3VX0
Xspi1_g932__5122 spi1_n_1929 spi1_Rx_count<4> spi1_n_1926 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg16857__2346 n_250 FE_PHN403_conf0_13 n_284 gnd3i! vdd3i! / NA2JI3VX0
Xg16856__2883 n_250 FE_PHN402_conf0_12 n_285 gnd3i! vdd3i! / NA2JI3VX0
Xg16859__7410 n_250 FE_PHN400_conf0_14 n_282 gnd3i! vdd3i! / NA2JI3VX0
Xg11868__1881 FE_OFN50_npg1_phase_up_state ele1<19> n_585 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11863__1705 npg1_phase_down_state ele2<19> n_590 gnd3i! vdd3i! / NA2JI3VX0
Xg11873__9315 npg1_phase_down_state ele2<18> n_580 gnd3i! vdd3i! / NA2JI3VX0
Xg11869__5115 FE_OFN50_npg1_phase_up_state ele1<18> n_584 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11880__5477 FE_OFN50_npg1_phase_up_state ele1<28> n_573 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11867__6131 npg1_phase_down_state ele2<28> n_586 gnd3i! vdd3i! / NA2JI3VX0
Xg11916__2883 FE_OFN50_npg1_phase_up_state ele1<17> n_551 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11878__7410 npg1_phase_down_state ele2<17> n_575 gnd3i! vdd3i! / NA2JI3VX0
Xg11921__5477 npg1_phase_down_state ele2<27> n_546 gnd3i! vdd3i! / NA2JI3VX0
Xg11917__2346 FE_OFN50_npg1_phase_up_state ele1<27> n_550 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11866__7098 npg1_phase_down_state ele2<26> n_587 gnd3i! vdd3i! / NA2JI3VX0
Xg11864__5122 FE_OFN50_npg1_phase_up_state ele1<26> n_589 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11877__1666 npg1_phase_down_state ele2<25> n_576 gnd3i! vdd3i! / NA2JI3VX0
Xg11872__6161 FE_OFN50_npg1_phase_up_state ele1<25> n_581 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11853__2398 FE_OFN57_npg1_phase_up_state ele2<2> n_600 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11854__5107 FE_OFN57_npg1_phase_up_state ele2<8> n_599 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11856__4319 FE_OFN57_npg1_phase_up_state ele2<6> n_597 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11857__8428 FE_OFN57_npg1_phase_up_state ele2<3> n_596 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11859__6783 FE_OFN50_npg1_phase_up_state ele2<17> n_594 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11860__3680 FE_OFN57_npg1_phase_up_state ele2<1> n_593 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11861__1617 FE_OFN57_npg1_phase_up_state ele2<9> n_592 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11862__2802 FE_OFN57_npg1_phase_up_state ele2<0> n_591 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11865__8246 FE_OFN50_npg1_phase_up_state ele2<19> n_588 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11871__4733 FE_OFN50_npg1_phase_up_state ele2<31> n_582 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11874__9945 FE_OFN50_npg1_phase_up_state ele2<21> n_579 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11879__6417 FE_OFN50_npg1_phase_up_state ele2<22> n_574 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11895__5107 FE_OFN57_npg1_phase_up_state ele2<7> n_572 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11898__8428 FE_OFN50_npg1_phase_up_state ele2<28> n_569 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11900__6783 FE_OFN50_npg1_phase_up_state ele2<23> n_567 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11901__3680 FE_OFN57_npg1_phase_up_state ele2<10> n_566 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11902__1617 FE_OFN50_npg1_phase_up_state ele2<18> n_565 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11903__2802 FE_OFN57_npg1_phase_up_state ele2<5> n_564 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11904__1705 FE_OFN57_npg1_phase_up_state ele2<11> n_563 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11905__5122 FE_OFN50_npg1_phase_up_state ele2<25> n_562 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11907__7098 FE_OFN50_npg1_phase_up_state ele2<24> n_560 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11908__6131 FE_OFN50_npg1_phase_up_state ele2<26> n_559 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11909__1881 FE_OFN50_npg1_phase_up_state ele2<30> n_558 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11911__7482 FE_OFN50_npg1_phase_up_state ele2<20> n_556 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11912__4733 FE_OFN50_npg1_phase_up_state ele2<27> n_555 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11913__6161 FE_OFN50_npg1_phase_up_state ele2<29> n_554 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11914__9315 FE_OFN57_npg1_phase_up_state ele2<4> n_553 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11915__9945 FE_OFN50_npg1_phase_up_state ele2<16> n_552 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11918__1666 FE_OFN57_npg1_phase_up_state ele2<12> n_549 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11919__7410 FE_OFN57_npg1_phase_up_state ele2<13> n_548 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11920__6417 FE_OFN57_npg1_phase_up_state ele2<14> n_547 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg11922__2398 FE_OFN50_npg1_phase_up_state ele2<15> n_545 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg16641__2802 n_443 npg1_OFF_count<9> n_463 gnd3i! vdd3i! / NA2JI3VX0
Xg16791__2398 n_10 npg1_DAC_cont<0> n_343 gnd3i! vdd3i! / NA2JI3VX0
Xg16643__5122 n_443 npg1_OFF_count<8> n_461 gnd3i! vdd3i! / NA2JI3VX0
Xg16733__1705 n_387 n_315 n_404 gnd3i! vdd3i! / NA2JI3VX0
Xg16942__8246 n_9 FE_OFN52_enable n_185 gnd3i! vdd3i! / NA2JI3VX0
Xg16955__1666 n_158 FE_OFN52_enable n_195 gnd3i! vdd3i! / NA2JI3VX0
Xg16991__6417 n_68 npg1_on_off_ctrl<1> n_160 gnd3i! vdd3i! / NA2JI3VX0
Xg16774__1881 n_347 npg1_OFF_count<7> n_361 gnd3i! vdd3i! / NA2JI3VX0
Xg16992__5477 n_69 npg1_OFF_count<2> n_159 gnd3i! vdd3i! / NA2JI3VX0
Xg17067__8428 n_34 conf0<25> n_85 gnd3i! vdd3i! / NA2JI3VX0
Xg16789__6417 n_10 npg1_DAC_cont<4> n_345 gnd3i! vdd3i! / NA2JI3VX0
Xg16790__5477 n_10 npg1_DAC_cont<3> n_344 gnd3i! vdd3i! / NA2JI3VX0
Xg16899__5107 n_225 n_40 n_237 gnd3i! vdd3i! / NA2JI3VX0
Xg16642__1705 n_444 npg1_ON_count<7> n_462 gnd3i! vdd3i! / NA2JI3VX0
Xg16809__7098 n_309 npg1_phase_up_count<2> n_325 gnd3i! vdd3i! / NA2JI3VX0
Xg16700__9945 n_406 FE_PHN399_npg1_freq_count_10 n_415 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg16667__7410 n_427 n_399 n_442 gnd3i! vdd3i! / NA2JI3VX0
Xg16654__8246 n_444 npg1_ON_count<6> n_459 gnd3i! vdd3i! / NA2JI3VX0
Xg16656__6131 n_447 npg1_ON_count<3> n_457 gnd3i! vdd3i! / NA2JI3VX0
Xg16831__2398 n_277 npg1_phase_up_count<1> n_307 gnd3i! vdd3i! / NA2JI3VX0
Xg16739__1881 n_371 npg1_freq_count<7> n_388 gnd3i! vdd3i! / NA2JI3VX0
Xg17038__1705 npg1_phase_up_count<2> n_56 n_108 gnd3i! vdd3i! / NA2JI3VX0
Xg17057__2883 npg1_freq_count<8> npg1_freq_count<7> n_59 gnd3i! vdd3i! / 
+ NA2JI3VX0
Xg16933__5526 n_204 npg1_ON_count<2> n_213 gnd3i! vdd3i! / NA2JI3VX0
Xg17075__8246 n_37 conf1<21> n_75 gnd3i! vdd3i! / NA2JI3VX0
Xg16923__2346 n_197 npg1_freq_count<4> n_222 gnd3i! vdd3i! / NA2JI3VX0
Xg16616__2883 n_460 npg1_UP_count<4> n_480 gnd3i! vdd3i! / NA2JI3VX0
Xg16633__5107 n_460 npg1_UP_count<5> n_473 gnd3i! vdd3i! / NA2JI3VX0
Xg16704__2346 n_324 n_407 n_424 gnd3i! vdd3i! / NA2JI3VX0
Xg16943__7098 n_160 FE_OFN52_enable n_184 gnd3i! vdd3i! / NA2JI3VX0
Xg16836__5526 n_275 FE_OFN52_enable n_312 gnd3i! vdd3i! / NA2JI3VX0
Xg16724__4319 n_396 npg1_DOWN_count<4> n_401 gnd3i! vdd3i! / NA2JI3VX0
Xg16725__8428 n_396 npg1_DOWN_count<5> n_400 gnd3i! vdd3i! / NA2JI3VX0
Xg17042__6131 n_18 conf0<2> n_103 gnd3i! vdd3i! / NA2JI3VX0
Xg16874__2802 n_267 npg1_UP_count<3> n_272 gnd3i! vdd3i! / NA2JI3VX0
Xg16873__1617 n_266 npg1_DOWN_count<3> n_273 gnd3i! vdd3i! / NA2JI3VX0
Xg17085__2883 npg1_UP_count<4> n_55 n_64 gnd3i! vdd3i! / NA2JI3VX0
Xg17084__9945 n_39 conf0<18> n_65 gnd3i! vdd3i! / NA2JI3VX0
Xg16801__3680 n_10 npg1_DAC_cont<5> n_333 gnd3i! vdd3i! / NA2JI3VX0
Xg16792__5107 n_10 npg1_DAC_cont<1> n_342 gnd3i! vdd3i! / NA2JI3VX0
Xg16793__6260 n_10 npg1_DAC_cont<2> n_341 gnd3i! vdd3i! / NA2JI3VX0
Xg16830__5477 n_279 npg1_phase_down_count<1> n_308 gnd3i! vdd3i! / NA2JI3VX0
Xg17062__5477 n_24 conf1<12> n_90 gnd3i! vdd3i! / NA2JI3VX0
Xg17059__1666 n_47 conf1<17> n_93 gnd3i! vdd3i! / NA2JI3VX0
Xg17063__2398 n_57 conf0<31> n_89 gnd3i! vdd3i! / NA2JI3VX0
Xg17073__1705 n_41 conf0<29> n_78 gnd3i! vdd3i! / NA2JI3VX0
Xg17060__7410 n_15 conf0<8> n_92 gnd3i! vdd3i! / NA2JI3VX0
Xg16917__7482 n_178 n_99 n_218 gnd3i! vdd3i! / NA2JI3VX0
Xg17078__1881 n_43 conf0<6> n_71 gnd3i! vdd3i! / NA2JI3VX0
Xg17089__7410 n_36 conf0<9> n_61 gnd3i! vdd3i! / NA2JI3VX0
Xg17045__5115 n_54 conf0<10> n_101 gnd3i! vdd3i! / NA2JI3VX0
Xg16637__5526 n_445 n_50 n_414 n_229 n_469 gnd3i! vdd3i! / ON22JI3VX1
Xg16999__6783 n_12 conf0<24> n_34 conf0<25> n_128 gnd3i! vdd3i! / ON22JI3VX1
Xg16638__6783 n_446 n_24 n_414 n_170 n_468 gnd3i! vdd3i! / ON22JI3VX1
Xg16745__9315 n_363 npg1_freq_count<8> n_15 npg1_freq_count<7> n_386 gnd3i! 
+ vdd3i! / ON22JI3VX1
Xg16752__5477 n_320 n_174 n_364 n_18 n_379 gnd3i! vdd3i! / ON22JI3VX1
Xg16751__6417 n_320 n_228 n_357 n_17 n_380 gnd3i! vdd3i! / ON22JI3VX1
Xg16819__4733 n_289 npg1_ON_count<4> n_16 npg1_ON_count<3> n_317 gnd3i! vdd3i! 
+ / ON22JI3VX1
Xg16844__1705 n_265 npg1_phase_up_count<0> n_37 n_66 n_299 gnd3i! vdd3i! / 
+ ON22JI3VX1
Xg16709__5477 n_394 n_36 n_393 npg1_freq_count<9> n_409 gnd3i! vdd3i! / 
+ ON22JI3VX1
Xg17008__1881 n_18 conf0<2> n_42 conf0<3> n_139 gnd3i! vdd3i! / ON22JI3VX1
Xg17005__8246 n_27 conf0<30> n_57 conf0<31> n_142 gnd3i! vdd3i! / ON22JI3VX1
Xg16869__8428 n_243 npg1_phase_down_count<0> npg1_phase_pause_ready 
+ FE_OFN58_npg1_phase_down_state n_279 gnd3i! vdd3i! / ON22JI3VX1
Xg17004__5122 n_48 conf1<16> n_47 conf1<17> n_143 gnd3i! vdd3i! / ON22JI3VX1
Xg17003__1705 n_43 conf0<6> n_38 conf0<7> n_144 gnd3i! vdd3i! / ON22JI3VX1
Xg16823__2883 n_271 n_270 n_102 n_160 n_321 gnd3i! vdd3i! / AN211JI3VX1
Xg16962__6260 npg1_UP_count<0> n_53 n_3 n_131 n_172 gnd3i! vdd3i! / AN211JI3VX1
Xg16949__4733 n_16 conf0<28> n_79 n_161 n_202 gnd3i! vdd3i! / AN211JI3VX1
Xg16970__2802 n_81 n_97 n_11 n_77 n_165 gnd3i! vdd3i! / AN211JI3VX1
Xg16971__1705 n_52 conf0<5> n_111 n_72 n_178 gnd3i! vdd3i! / AN211JI3VX1
Xspi1_g993 spi1_Rx_count<0> spi1_n_2088 gnd3i! vdd3i! / INJI3VX0
Xg11954 ele1<2> n_514 gnd3i! vdd3i! / INJI3VX0
Xg11932 ele1<8> n_536 gnd3i! vdd3i! / INJI3VX0
Xg11946 ele1<6> n_522 gnd3i! vdd3i! / INJI3VX0
Xg11948 ele1<3> n_520 gnd3i! vdd3i! / INJI3VX0
Xg11928 ele1<17> n_540 gnd3i! vdd3i! / INJI3VX0
Xg11933 ele1<1> n_535 gnd3i! vdd3i! / INJI3VX0
Xg11942 ele1<9> n_526 gnd3i! vdd3i! / INJI3VX0
Xg11938 ele1<0> n_530 gnd3i! vdd3i! / INJI3VX0
Xg11925 ele1<19> n_543 gnd3i! vdd3i! / INJI3VX0
Xg11934 ele1<31> n_534 gnd3i! vdd3i! / INJI3VX0
Xg11936 ele1<21> n_532 gnd3i! vdd3i! / INJI3VX0
Xg11939 ele1<22> n_529 gnd3i! vdd3i! / INJI3VX0
Xg11950 ele1<7> n_518 gnd3i! vdd3i! / INJI3VX0
Xg11951 ele1<28> n_517 gnd3i! vdd3i! / INJI3VX0
Xg11953 ele1<23> n_515 gnd3i! vdd3i! / INJI3VX0
Xg11952 ele1<10> n_516 gnd3i! vdd3i! / INJI3VX0
Xg11945 ele1<18> n_523 gnd3i! vdd3i! / INJI3VX0
Xg11947 ele1<5> n_521 gnd3i! vdd3i! / INJI3VX0
Xg11943 ele1<11> n_525 gnd3i! vdd3i! / INJI3VX0
Xg11929 ele1<25> n_539 gnd3i! vdd3i! / INJI3VX0
Xg11940 ele1<24> n_528 gnd3i! vdd3i! / INJI3VX0
Xg11927 ele1<26> n_541 gnd3i! vdd3i! / INJI3VX0
Xg11949 ele1<30> n_519 gnd3i! vdd3i! / INJI3VX0
Xg11930 ele1<20> n_538 gnd3i! vdd3i! / INJI3VX0
Xg11944 ele1<27> n_524 gnd3i! vdd3i! / INJI3VX0
Xg11935 ele1<29> n_533 gnd3i! vdd3i! / INJI3VX0
Xg11926 ele1<4> n_542 gnd3i! vdd3i! / INJI3VX0
Xg11955 ele1<16> n_513 gnd3i! vdd3i! / INJI3VX0
Xg11937 ele1<12> n_531 gnd3i! vdd3i! / INJI3VX0
Xg11924 ele1<13> n_544 gnd3i! vdd3i! / INJI3VX0
Xg11931 ele1<14> n_537 gnd3i! vdd3i! / INJI3VX0
Xg11941 ele1<15> n_527 gnd3i! vdd3i! / INJI3VX0
Xg16734 n_361 n_397 gnd3i! vdd3i! / INJI3VX0
Xg16887 n_250 n_249 gnd3i! vdd3i! / INJI3VX0
Xg16972 n_6 n_164 gnd3i! vdd3i! / INJI3VX0
Xg16877 n_262 n_261 gnd3i! vdd3i! / INJI3VX0
Xg16705 n_414 n_413 gnd3i! vdd3i! / INJI3VX0
Xg16722 n_404 n_403 gnd3i! vdd3i! / INJI3VX0
Xg17101 npg1_OFF_count<4> n_50 gnd3i! vdd3i! / INJI3VX0
Xg17102 npg1_OFF_count<1> n_49 gnd3i! vdd3i! / INJI3VX0
Xg17129 npg1_OFF_count<2> n_24 gnd3i! vdd3i! / INJI3VX0
Xg16694 n_426 n_425 gnd3i! vdd3i! / INJI3VX0
Xg17119 npg1_ON_count<1> n_34 gnd3i! vdd3i! / INJI3VX0
Xg17147 npg1_ON_count<0> n_12 gnd3i! vdd3i! / INJI3VX0
Xg17128 npg1_DOWN_accumulator<4> n_25 gnd3i! vdd3i! / INJI3VX0
Xg17112 npg1_phase_pause_ready n_40 gnd3i! vdd3i! / INJI3VX0
Xg16912 n_225 n_226 gnd3i! vdd3i! / INJI3VX0
Xg16863 n_277 n_278 gnd3i! vdd3i! / INJI3VX0
Xg16768 n_362 n_363 gnd3i! vdd3i! / INJI3VX0
Xg17144 npg1_freq_count<8> n_15 gnd3i! vdd3i! / INJI3VX0
Xg17140 npg1_freq_count<2> n_18 gnd3i! vdd3i! / INJI3VX0
Xg16864 n_275 n_276 gnd3i! vdd3i! / INJI3VX0
Xg17091 conf1<23> n_56 gnd3i! vdd3i! / INJI3VX0
Xg17124 npg1_phase_up_count<2> n_29 gnd3i! vdd3i! / INJI3VX0
Xg17114 npg1_freq_count<7> n_38 gnd3i! vdd3i! / INJI3VX0
Xg16767 n_365 n_366 gnd3i! vdd3i! / INJI3VX0
Xg17143 npg1_ON_count<4> n_16 gnd3i! vdd3i! / INJI3VX0
Xg17115 npg1_phase_up_count<0> n_37 gnd3i! vdd3i! / INJI3VX0
Xg17100 npg1_phase_up_count<1> n_51 gnd3i! vdd3i! / INJI3VX0
Xg16817 n_320 n_319 gnd3i! vdd3i! / INJI3VX0
Xg17118 npg1_freq_count<1> n_35 gnd3i! vdd3i! / INJI3VX0
Xg17117 npg1_freq_count<9> n_36 gnd3i! vdd3i! / INJI3VX0
Xg16805 n_272 n_331 gnd3i! vdd3i! / INJI3VX0
Xg17127 conf0<19> n_26 gnd3i! vdd3i! / INJI3VX0
Xg17145 npg1_DOWN_count<4> n_14 gnd3i! vdd3i! / INJI3VX0
Xg17120 npg1_UP_count<0> n_33 gnd3i! vdd3i! / INJI3VX0
Xg17095 conf0<18> n_53 gnd3i! vdd3i! / INJI3VX0
Xg17015 n_104 n_105 gnd3i! vdd3i! / INJI3VX0
Xg17017 n_5 n_98 gnd3i! vdd3i! / INJI3VX0
Xg16806 n_273 n_330 gnd3i! vdd3i! / INJI3VX0
Xg16688 n_431 n_430 gnd3i! vdd3i! / INJI3VX0
Xg16695 n_424 n_423 gnd3i! vdd3i! / INJI3VX0
Xg16796 n_339 n_338 gnd3i! vdd3i! / INJI3VX0
Xg17093 conf0<22> n_55 gnd3i! vdd3i! / INJI3VX0
Xg16778 n_356 n_355 gnd3i! vdd3i! / INJI3VX0
Xg17113 npg1_DOWN_count<0> n_39 gnd3i! vdd3i! / INJI3VX0
Xg17130 npg1_DOWN_count<2> n_23 gnd3i! vdd3i! / INJI3VX0
Xg17132 npg1_DOWN_count<1> n_21 gnd3i! vdd3i! / INJI3VX0
Xg17146 npg1_freq_count<0> n_13 gnd3i! vdd3i! / INJI3VX0
Xg17142 npg1_freq_count<4> n_17 gnd3i! vdd3i! / INJI3VX0
Xg17122 conf0<16> n_31 gnd3i! vdd3i! / INJI3VX0
Xg17123 conf0<15> n_30 gnd3i! vdd3i! / INJI3VX0
Xg16875 n_235 n_268 gnd3i! vdd3i! / INJI3VX0
Xg16934 n_96 n_203 gnd3i! vdd3i! / INJI3VX0
Xg16935 n_200 n_201 gnd3i! vdd3i! / INJI3VX0
Xg16973 n_161 n_162 gnd3i! vdd3i! / INJI3VX0
Xg17053 n_78 n_79 gnd3i! vdd3i! / INJI3VX0
Xg17125 npg1_phase_down_count<2> n_28 gnd3i! vdd3i! / INJI3VX0
Xg17051 n_93 n_94 gnd3i! vdd3i! / INJI3VX0
Xg16876 n_264 n_263 gnd3i! vdd3i! / INJI3VX0
Xg17105 npg1_OFF_count<5> n_46 gnd3i! vdd3i! / INJI3VX0
Xg17103 npg1_OFF_count<6> n_48 gnd3i! vdd3i! / INJI3VX0
Xg17104 npg1_OFF_count<7> n_47 gnd3i! vdd3i! / INJI3VX0
Xg17090 npg1_ON_count<7> n_57 gnd3i! vdd3i! / INJI3VX0
Xg17126 npg1_ON_count<6> n_27 gnd3i! vdd3i! / INJI3VX0
Xg17111 npg1_ON_count<5> n_41 gnd3i! vdd3i! / INJI3VX0
Xg17107 npg1_phase_down_count<0> n_45 gnd3i! vdd3i! / INJI3VX0
Xg17054 n_76 n_77 gnd3i! vdd3i! / INJI3VX0
Xg17055 n_71 n_72 gnd3i! vdd3i! / INJI3VX0
Xg16798__8428 n_300 n_11 n_249 n_195 n_336 gnd3i! vdd3i! / ON211JI3VX1
Xg16832__5107 n_242 n_195 n_274 n_220 n_306 gnd3i! vdd3i! / ON211JI3VX1
Xg16852__4733 n_6 FE_OFN52_enable n_249 n_261 n_291 gnd3i! vdd3i! / ON211JI3VX1
Xg16754__5107 n_358 n_121 n_134 n_87 n_387 gnd3i! vdd3i! / ON211JI3VX1
Xg16728__3680 n_368 n_119 n_158 n_88 n_407 gnd3i! vdd3i! / ON211JI3VX1
Xg16957__7410 n_39 conf0<18> n_148 n_113 n_177 gnd3i! vdd3i! / ON211JI3VX1
Xg16947__5115 n_13 conf0<0> n_105 n_103 n_181 gnd3i! vdd3i! / ON211JI3VX1
Xg16928__2398 n_62 n_65 n_138 n_5 n_208 gnd3i! vdd3i! / ON211JI3VX1
Xg16897__5477 n_113 n_98 n_208 n_122 n_245 gnd3i! vdd3i! / ON211JI3VX1
Xg16635__4319 n_433 n_263 n_333 n_294 n_471 gnd3i! vdd3i! / ON211JI3VX1
Xg16658__5115 n_418 n_263 n_345 n_295 n_455 gnd3i! vdd3i! / ON211JI3VX1
Xg16707__7410 n_263 n_377 n_344 n_296 n_411 gnd3i! vdd3i! / ON211JI3VX1
Xg16994__5107 n_22 conf1<22> n_45 conf1<21> n_133 gnd3i! vdd3i! / ON211JI3VX1
Xg16926__6417 n_67 n_104 n_163 n_61 n_210 gnd3i! vdd3i! / ON211JI3VX1
Xg16858__1666 n_186 n_111 n_247 n_218 n_283 gnd3i! vdd3i! / ON211JI3VX1
Xg16699__9315 n_397 npg1_OFF_count<8> npg1_OFF_count<9> n_416 gnd3i! vdd3i! / 
+ AN21JI3VX1
Xg16671__5107 n_413 n_159 n_403 n_445 gnd3i! vdd3i! / AN21JI3VX1
Xg16741__7482 n_359 n_231 n_9 n_395 gnd3i! vdd3i! / AN21JI3VX1
Xg16812__5115 n_280 n_123 n_110 n_322 gnd3i! vdd3i! / AN21JI3VX1
Xg16976__7098 n_12 conf0<24> n_100 n_155 gnd3i! vdd3i! / AN21JI3VX1
Xg16843__2802 n_252 n_134 n_164 n_300 gnd3i! vdd3i! / AN21JI3VX1
Xg16732__2802 n_312 n_185 n_395 n_405 gnd3i! vdd3i! / AN21JI3VX1
Xg16737__7098 n_365 npg1_ON_count<6> npg1_ON_count<7> n_390 gnd3i! vdd3i! / 
+ AN21JI3VX1
Xg16786__2346 n_319 n_135 n_11 n_357 gnd3i! vdd3i! / AN21JI3VX1
Xg16884__5115 n_739 FE_OFN50_npg1_phase_up_state npg1_pulse_start n_265 gnd3i! 
+ vdd3i! / AN21JI3VX1
Xg16742__4733 n_319 n_59 n_371 n_394 gnd3i! vdd3i! / AN21JI3VX1
Xg16780__7482 n_331 npg1_UP_count<4> npg1_UP_count<5> n_353 gnd3i! vdd3i! / 
+ AN21JI3VX1
Xg16868__4319 n_239 n_4 n_205 n_269 gnd3i! vdd3i! / AN21JI3VX1
Xg16804__1705 n_312 n_184 n_321 n_339 gnd3i! vdd3i! / AN21JI3VX1
Xg16866__5107 n_245 npg1_DOWN_count<4> n_109 n_271 gnd3i! vdd3i! / AN21JI3VX1
Xg16995__6260 n_33 conf0<18> n_63 n_132 gnd3i! vdd3i! / AN21JI3VX1
Xg16782__6161 n_330 npg1_DOWN_count<4> npg1_DOWN_count<5> n_351 gnd3i! vdd3i! 
+ / AN21JI3VX1
Xg17171 n_17 conf0<4> n_743 n_744 gnd3i! vdd3i! / AN21JI3VX1
Xg16853__6161 n_268 n_115 n_82 n_290 gnd3i! vdd3i! / AN21JI3VX1
Xg16911__7098 n_80 n_203 n_116 n_235 gnd3i! vdd3i! / AN21JI3VX1
Xg16888__6161 n_206 n_86 n_112 n_248 gnd3i! vdd3i! / AN21JI3VX1
Xg16896__6417 n_201 n_107 n_212 n_238 gnd3i! vdd3i! / AN21JI3VX1
Xg16931__4319 n_50 conf1<14> n_200 n_215 gnd3i! vdd3i! / AN21JI3VX1
Xg17006__7098 n_48 conf1<16> n_94 n_141 gnd3i! vdd3i! / AN21JI3VX1
Xg16892__2346 n_214 FE_OFN58_npg1_phase_down_state npg1_phase_pause_ready 
+ n_251 gnd3i! vdd3i! / AN21JI3VX1
Xg16941__5122 n_71 n_74 n_144 n_186 gnd3i! vdd3i! / AN21JI3VX1
Xspi1_g987__9945 spi1_Rx_count<2> spi1_Rx_count<3> spi1_n_2017 spi1_n_2010 
+ gnd3i! vdd3i! / NA3I1JI3VX1
Xg17168 FE_OFN58_npg1_phase_down_state n_40 npg1_phase_down_count<0> n_740 
+ gnd3i! vdd3i! / NA3I1JI3VX1
Xg16965__5526 n_70 n_85 n_155 n_169 gnd3i! vdd3i! / NA3I1JI3VX1
Xg17001__1617 npg1_phase_up_count<2> npg1_phase_up_count<0> 
+ npg1_phase_up_count<1> n_126 gnd3i! vdd3i! / NA3I1JI3VX1
Xg16726__5526 n_393 npg1_freq_count<9> FE_PHN399_npg1_freq_count_10 n_399 
+ gnd3i! vdd3i! / NA3I1JI3VX1
Xg16871__6783 n_7 n_232 n_233 n_275 gnd3i! vdd3i! / NA3I1JI3VX1
Xg16959__5477 n_106 n_92 n_137 n_175 gnd3i! vdd3i! / NA3I1JI3VX1
Xg17000__3680 npg1_phase_down_count<2> npg1_phase_down_count<0> 
+ npg1_phase_down_count<1> n_127 gnd3i! vdd3i! / NA3I1JI3VX1
Xg17151__5107 n_81 n_101 n_151 n_7 gnd3i! vdd3i! / NA3I1JI3VX1
Xg16784__9945 n_285 n_297 n_343 n_349 gnd3i! vdd3i! / NA3JI3VX0
Xg16690__7098 FE_PHN405_npg1_OFF_count_0 n_49 n_413 n_428 gnd3i! vdd3i! / 
+ NA3JI3VX0
Xg16711__5107 n_404 n_387 FE_OFN52_enable n_414 gnd3i! vdd3i! / NA3JI3VX0
Xg16799__5526 npg1_freq_count<0> n_35 n_319 n_335 gnd3i! vdd3i! / NA3JI3VX0
Xg17012__6161 npg1_freq_count<2> npg1_freq_count<1> npg1_freq_count<0> n_135 
+ gnd3i! vdd3i! / NA3JI3VX0
Xg16743__6161 npg1_freq_count<8> n_362 n_319 n_393 gnd3i! vdd3i! / NA3JI3VX0
Xg16958__6417 n_122 n_5 n_138 n_176 gnd3i! vdd3i! / NA3JI3VX0
Xg16966__6783 n_64 n_0 n_132 n_168 gnd3i! vdd3i! / NA3JI3VX0
Xg16693__5115 FE_OFN52_enable n_407 n_424 n_431 gnd3i! vdd3i! / NA3JI3VX0
Xg16783__9315 n_284 n_298 n_342 n_350 gnd3i! vdd3i! / NA3JI3VX0
Xg16736__8246 n_282 n_348 n_341 n_391 gnd3i! vdd3i! / NA3JI3VX0
Xg16914__6131 n_136 n_149 n_173 n_221 gnd3i! vdd3i! / NA3JI3VX0
Xg16969__1617 n_76 n_97 n_150 n_166 gnd3i! vdd3i! / NA3JI3VX0
Xg16825__2346 n_311 n_210 n_165 n_320 gnd3i! vdd3i! / NA3JI3VX0
Xspi1_g940__5115 spi1_n_1998 spi1_Rx_data_temp<32> spi1_n_1995 gnd3i! vdd3i! / 
+ NO2I1JI3VX1
Xg16974__5122 n_85 conf0<24> n_157 gnd3i! vdd3i! / NO2I1JI3VX1
Xg16886__4733 n_242 n_195 n_262 gnd3i! vdd3i! / NO2I1JI3VX1
Xg16885__7482 n_236 n_196 n_264 gnd3i! vdd3i! / NO2I1JI3VX1
Xg17022__7410 npg1_OFF_count<9> conf1<19> n_121 gnd3i! vdd3i! / NO2I1JI3VX1
Xg17157__3680 npg1_ON_count<3> conf0<27> n_1 gnd3i! vdd3i! / NO2I1JI3VX1
Xg17035__1617 conf0<27> npg1_ON_count<3> n_110 gnd3i! vdd3i! / NO2I1JI3VX1
Xg17019__2883 conf0<20> npg1_UP_count<2> n_124 gnd3i! vdd3i! / NO2I1JI3VX1
Xg17024__5477 npg1_UP_count<5> conf0<23> n_119 gnd3i! vdd3i! / NO2I1JI3VX1
Xg17037__2802 npg1_DOWN_count<5> conf0<23> n_109 gnd3i! vdd3i! / NO2I1JI3VX1
Xg17043__1881 conf0<23> npg1_DOWN_count<5> n_102 gnd3i! vdd3i! / NO2I1JI3VX1
Xg16983__9315 n_65 n_62 n_148 gnd3i! vdd3i! / NO2I1JI3VX1
Xg17155__5526 npg1_UP_count<2> conf0<20> n_3 gnd3i! vdd3i! / NO2I1JI3VX1
Xg16982__6161 n_90 n_117 n_149 gnd3i! vdd3i! / NO2I1JI3VX1
Xg17027__6260 conf0<13> npg1_DOWN_accumulator<5> n_116 gnd3i! vdd3i! / 
+ NO2I1JI3VX1
Xg17070__3680 conf0<14> npg1_DOWN_accumulator<6> n_82 gnd3i! vdd3i! / 
+ NO2I1JI3VX1
Xg17061__6417 conf1<18> npg1_OFF_count<8> n_91 gnd3i! vdd3i! / NO2I1JI3VX1
Xg16981__4733 n_61 n_67 n_150 gnd3i! vdd3i! / NO2I1JI3VX1
Xg11744__2802 n_635 n_637 n_634 n_636 n_644 gnd3i! vdd3i! / NA4JI3VX0
Xg16920__9315 n_140 n_108 n_75 n_153 n_225 gnd3i! vdd3i! / NA4JI3VX0
Xg16901__4319 n_172 n_88 n_120 n_207 n_242 gnd3i! vdd3i! / NA4JI3VX0
Xg16826__1666 n_163 n_92 n_61 n_283 n_311 gnd3i! vdd3i! / NA4JI3VX0
Xg17166 n_214 FE_OFN58_npg1_phase_down_state n_40 n_738 gnd3i! vdd3i! / 
+ NA22JI3VX1
Xg16673__4319 n_361 n_413 n_404 n_443 gnd3i! vdd3i! / NA22JI3VX1
Xg16766__2802 n_313 n_319 enable n_371 gnd3i! vdd3i! / NA22JI3VX1
Xg17172 n_42 conf0<3> n_178 n_743 gnd3i! vdd3i! / NA22JI3VX1
Xg16666__1666 n_272 n_430 n_424 n_460 gnd3i! vdd3i! / NA22JI3VX1
Xg16740__5115 n_273 n_356 n_338 n_396 gnd3i! vdd3i! / NA22JI3VX1
Xg16950__6161 conf1<15> n_46 n_141 n_200 gnd3i! vdd3i! / NA22JI3VX1
Xg16988__1666 conf0<30> n_27 n_89 n_161 gnd3i! vdd3i! / NA22JI3VX1
Xg16655__7098 n_445 FE_PHN397_npg1_OFF_count_3 n_458 gnd3i! vdd3i! / 
+ NA2I1JI3VX1
Xg16763__6783 n_357 FE_PHN398_npg1_freq_count_3 n_369 gnd3i! vdd3i! / 
+ NA2I1JI3VX1
Xg16979__5115 n_121 n_87 n_152 gnd3i! vdd3i! / NA2I1JI3VX1
Xg17065__6260 npg1_OFF_count<9> conf1<19> n_87 gnd3i! vdd3i! / NA2I1JI3VX1
Xg17020__2346 conf0<26> npg1_ON_count<2> n_123 gnd3i! vdd3i! / NA2I1JI3VX1
Xg17156__6783 npg1_ON_count<2> conf0<26> n_2 gnd3i! vdd3i! / NA2I1JI3VX1
Xg17149__5477 n_114 npg1_on_off_ctrl<1> n_9 gnd3i! vdd3i! / NA2I1JI3VX1
Xg17029__8428 npg1_on_off_ctrl<2> npg1_on_off_ctrl<0> n_114 gnd3i! vdd3i! / 
+ NA2I1JI3VX1
Xg17152__6260 npg1_on_off_ctrl<1> n_68 n_6 gnd3i! vdd3i! / NA2I1JI3VX1
Xg16862__2398 n_213 npg1_ON_count<3> n_289 gnd3i! vdd3i! / NA2I1JI3VX1
Xg17021__1666 conf0<21> npg1_DOWN_count<3> n_122 gnd3i! vdd3i! / NA2I1JI3VX1
Xg17023__6417 conf0<21> npg1_UP_count<3> n_120 gnd3i! vdd3i! / NA2I1JI3VX1
Xg17049__6161 npg1_freq_count<11> conf0<11> n_97 gnd3i! vdd3i! / NA2I1JI3VX1
Xg16834__4319 n_241 npg1_freq_count<6> n_313 gnd3i! vdd3i! / NA2I1JI3VX1
Xg16902__8428 n_222 npg1_freq_count<5> n_241 gnd3i! vdd3i! / NA2I1JI3VX1
Xg17064__5107 npg1_UP_count<5> conf0<23> n_88 gnd3i! vdd3i! / NA2I1JI3VX1
Xg17154__8428 npg1_UP_count<1> conf0<19> n_4 gnd3i! vdd3i! / NA2I1JI3VX1
Xg17158__1617 npg1_UP_count<3> conf0<21> n_0 gnd3i! vdd3i! / NA2I1JI3VX1
Xg17153__4319 npg1_DOWN_count<3> conf0<21> n_5 gnd3i! vdd3i! / NA2I1JI3VX1
Xg17074__5122 conf0<11> npg1_freq_count<11> n_76 gnd3i! vdd3i! / NA2I1JI3VX1
Xg16989__7410 n_82 n_115 n_145 gnd3i! vdd3i! / NA2I1JI3VX1
Xg16987__2346 n_116 n_80 n_146 gnd3i! vdd3i! / NA2I1JI3VX1
Xg16984__9945 n_91 n_73 n_147 gnd3i! vdd3i! / NA2I1JI3VX1
Xg17072__2802 conf0<13> npg1_DOWN_accumulator<5> n_80 gnd3i! vdd3i! / 
+ NA2I1JI3VX1
Xg17028__4319 conf0<14> npg1_DOWN_accumulator<6> n_115 gnd3i! vdd3i! / 
+ NA2I1JI3VX1
Xg17077__6131 conf1<18> npg1_OFF_count<8> n_73 gnd3i! vdd3i! / NA2I1JI3VX1
Xg16954__2346 n_160 n_11 n_196 gnd3i! vdd3i! / OR2JI3VX0
Xg16951__9315 n_9 n_11 n_199 gnd3i! vdd3i! / OR2JI3VX0
Xg17083__9315 FE_OFN50_npg1_phase_up_state npg1_pulse_start n_66 gnd3i! vdd3i! 
+ / OR2JI3VX0
Xg17030__5526 n_23 conf0<20> n_113 gnd3i! vdd3i! / OR2JI3VX0
Xg17066__4319 n_24 conf1<12> n_86 gnd3i! vdd3i! / OR2JI3VX0
XFE_OFC76_DAC_3 FE_OFN45_DAC_3 DAC<3> gnd3i! vdd3i! / BUJI3VX12
XFE_OFC75_DAC_2 FE_OFN44_DAC_2 DAC<2> gnd3i! vdd3i! / BUJI3VX12
XFE_OFC74_DAC_1 FE_OFN43_DAC_1 DAC<1> gnd3i! vdd3i! / BUJI3VX12
Xg11739__5526 FE_OFN39_pulse_active npg1_DAC_cont<0> FE_OFN42_DAC_0 gnd3i! 
+ vdd3i! / AND2JI3VX1
Xg11735__5107 FE_OFN39_pulse_active npg1_DAC_cont<4> FE_OFN46_DAC_4 gnd3i! 
+ vdd3i! / AND2JI3VX1
Xg11734__2398 FE_OFN39_pulse_active npg1_DAC_cont<5> FE_OFN47_DAC_5 gnd3i! 
+ vdd3i! / AND2JI3VX1
Xg11736__6260 FE_OFN39_pulse_active npg1_DAC_cont<3> FE_OFN45_DAC_3 gnd3i! 
+ vdd3i! / AND2JI3VX1
Xg11737__4319 FE_OFN39_pulse_active npg1_DAC_cont<2> FE_OFN44_DAC_2 gnd3i! 
+ vdd3i! / AND2JI3VX1
Xg11738__8428 FE_OFN39_pulse_active npg1_DAC_cont<1> FE_OFN43_DAC_1 gnd3i! 
+ vdd3i! / AND2JI3VX1
XFE_PHC432_n_32 FE_PHN422_n_32 FE_PHN432_n_32 gnd3i! vdd3i! / BUJI3VX8
XFE_PHC437_n_32 FE_PHN422_n_32 FE_PHN437_n_32 gnd3i! vdd3i! / BUJI3VX8
XCTS_ccl_a_buf_00004 CTS_3 CTS_2 gnd3i! vdd3i! / BUJI3VX8
XCTS_ccl_a_buf_00003 CTS_3 CTS_1 gnd3i! vdd3i! / BUJI3VX8
XCTS_ccl_a_buf_00002 CTS_3 CTS_5 gnd3i! vdd3i! / BUJI3VX8
XCTS_ccl_a_buf_00001 CTS_3 CTS_4 gnd3i! vdd3i! / BUJI3VX8
XFE_OFC98_OFN42_DAC_0 FE_OFN42_DAC_0 DAC<0> gnd3i! vdd3i! / BUJI3VX8
XFE_OFC97_OFN46_DAC_4 FE_OFN46_DAC_4 DAC<4> gnd3i! vdd3i! / BUJI3VX8
XFE_OFC96_OFN47_DAC_5 FE_OFN47_DAC_5 DAC<5> gnd3i! vdd3i! / BUJI3VX8
Xg16861__5477 n_204 n_219 n_157 n_2 n_280 gnd3i! vdd3i! / ON31JI3VX1
Xg16631__5477 npg1_OFF_count<8> n_361 n_414 n_461 n_475 gnd3i! vdd3i! / 
+ ON31JI3VX1
Xg16630__6417 npg1_OFF_count<3> n_159 n_414 n_458 n_476 gnd3i! vdd3i! / 
+ ON31JI3VX1
Xg16689__8246 npg1_freq_count<10> n_36 n_393 n_415 n_429 gnd3i! vdd3i! / 
+ ON31JI3VX1
Xg16632__2398 npg1_ON_count<6> n_366 n_425 n_459 n_474 gnd3i! vdd3i! / 
+ ON31JI3VX1
Xg16628__1666 npg1_ON_count<3> n_213 n_425 n_457 n_478 gnd3i! vdd3i! / 
+ ON31JI3VX1
Xg16822__9945 npg1_phase_up_count<1> n_37 n_265 n_307 n_314 gnd3i! vdd3i! / 
+ ON31JI3VX1
Xg16727__6783 npg1_freq_count<7> n_313 n_320 n_388 n_398 gnd3i! vdd3i! / 
+ ON31JI3VX1
Xg16738__6131 npg1_freq_count<3> n_135 n_320 n_369 n_389 gnd3i! vdd3i! / 
+ ON31JI3VX1
Xg16608__4733 npg1_UP_count<4> n_272 n_431 n_480 n_484 gnd3i! vdd3i! / 
+ ON31JI3VX1
Xg16706__1666 npg1_DOWN_count<4> n_273 n_355 n_401 n_412 gnd3i! vdd3i! / 
+ ON31JI3VX1
Xg16818__7482 npg1_phase_down_count<1> n_45 n_251 n_308 n_318 gnd3i! vdd3i! / 
+ ON31JI3VX1
Xg11845__2883 n_510 ele2<22> FE_OFN50_npg1_phase_up_state ele1<22> n_607 
+ gnd3i! vdd3i! / AN22JI3VX1
Xg11808__2883 n_509 ele2<15> FE_OFN50_npg1_phase_up_state ele1<15> n_612 
+ gnd3i! vdd3i! / AN22JI3VX1
Xg11849__6417 n_509 ele2<14> FE_OFN57_npg1_phase_up_state ele1<14> n_603 
+ gnd3i! vdd3i! / AN22JI3VX1
Xg16908__1705 n_198 n_50 npg1_OFF_count<4> FE_PHN233_npg1_OFF_count_3 n_229 
+ gnd3i! vdd3i! / AN22JI3VX1
Xg16846__8246 n_264 n_156 n_262 npg1_UP_accumulator<4> n_297 gnd3i! vdd3i! / 
+ AN22JI3VX1
Xg16964__8428 n_69 n_24 n_49 npg1_OFF_count<2> n_170 gnd3i! vdd3i! / AN22JI3VX1
Xg16960__2398 n_60 npg1_freq_count<0> n_35 npg1_freq_count<2> n_174 gnd3i! 
+ vdd3i! / AN22JI3VX1
Xg16909__5122 n_197 n_17 n_42 npg1_freq_count<4> n_228 gnd3i! vdd3i! / 
+ AN22JI3VX1
Xg17007__6131 n_29 conf1<23> n_51 conf1<22> n_140 gnd3i! vdd3i! / AN22JI3VX1
Xg17002__2802 npg1_DOWN_count<4> n_55 n_14 conf0<22> n_125 gnd3i! vdd3i! / 
+ AN22JI3VX1
Xg17010__7482 n_35 conf0<1> n_13 conf0<0> n_137 gnd3i! vdd3i! / AN22JI3VX1
Xg17009__5115 n_23 conf0<20> n_21 conf0<19> n_138 gnd3i! vdd3i! / AN22JI3VX1
Xg16849__1881 n_250 conf0<17> n_262 npg1_UP_accumulator<9> n_294 gnd3i! vdd3i! 
+ / AN22JI3VX1
Xg16845__5122 n_264 n_234 n_262 npg1_UP_accumulator<5> n_298 gnd3i! vdd3i! / 
+ AN22JI3VX1
Xg16785__2883 n_264 n_303 n_262 npg1_UP_accumulator<6> n_348 gnd3i! vdd3i! / 
+ AN22JI3VX1
Xg16848__6131 n_250 conf0<16> n_262 npg1_UP_accumulator<8> n_295 gnd3i! vdd3i! 
+ / AN22JI3VX1
Xg16847__7098 n_250 conf0<15> n_262 npg1_UP_accumulator<7> n_296 gnd3i! vdd3i! 
+ / AN22JI3VX1
Xg17011__4733 n_49 conf1<11> n_44 conf1<10> n_136 gnd3i! vdd3i! / AN22JI3VX1
Xg16906__1617 n_162 n_8 n_142 n_89 n_231 gnd3i! vdd3i! / AN22JI3VX1
Xg16932__8428 n_130 n_133 npg1_phase_down_count<2> n_56 n_214 gnd3i! vdd3i! / 
+ AN22JI3VX1
Xg16997__8428 n_28 conf1<23> n_22 conf1<22> n_130 gnd3i! vdd3i! / AN22JI3VX1
Xg11794__1617 n_590 FE_OFN50_npg1_phase_up_state n_585 FE_OFN12_up_switches_19 
+ gnd3i! vdd3i! / ON21JI3VX1
Xg11804__4733 n_580 FE_OFN50_npg1_phase_up_state n_584 FE_OFN13_up_switches_18 
+ gnd3i! vdd3i! / ON21JI3VX1
Xg11806__9315 n_586 FE_OFN50_npg1_phase_up_state n_573 FE_OFN4_up_switches_28 
+ gnd3i! vdd3i! / ON21JI3VX1
Xg11807__9945 n_575 FE_OFN50_npg1_phase_up_state n_551 FE_OFN14_up_switches_17 
+ gnd3i! vdd3i! / ON21JI3VX1
Xg16842__1617 n_251 npg1_phase_down_count<0> n_740 n_301 gnd3i! vdd3i! / 
+ ON21JI3VX1
Xg11788__6260 n_546 FE_OFN50_npg1_phase_up_state n_550 FE_OFN5_up_switches_27 
+ gnd3i! vdd3i! / ON21JI3VX1
Xg11790__8428 n_587 FE_OFN50_npg1_phase_up_state n_589 FE_OFN6_up_switches_26 
+ gnd3i! vdd3i! / ON21JI3VX1
Xg11795__2802 n_576 FE_OFN50_npg1_phase_up_state n_581 FE_OFN7_up_switches_25 
+ gnd3i! vdd3i! / ON21JI3VX1
Xg16627__2346 n_414 n_416 n_463 n_479 gnd3i! vdd3i! / ON21JI3VX1
Xg16770__5122 n_322 n_1 n_202 n_359 gnd3i! vdd3i! / ON21JI3VX1
Xg16629__7410 n_446 n_49 n_428 n_477 gnd3i! vdd3i! / ON21JI3VX1
Xg16821__9315 n_134 n_11 n_312 n_315 gnd3i! vdd3i! / ON21JI3VX1
Xg16841__3680 n_236 n_196 n_274 n_302 gnd3i! vdd3i! / ON21JI3VX1
Xg16634__6260 n_425 n_390 n_462 n_472 gnd3i! vdd3i! / ON21JI3VX1
Xg16829__6417 n_244 npg1_phase_up_count<1> n_278 n_309 gnd3i! vdd3i! / 
+ ON21JI3VX1
Xg16802__1617 n_265 n_126 n_325 n_332 gnd3i! vdd3i! / ON21JI3VX1
Xg16691__6131 n_406 n_319 npg1_freq_count<11> n_427 gnd3i! vdd3i! / ON21JI3VX1
Xg16735__5122 n_364 n_35 n_335 n_392 gnd3i! vdd3i! / ON21JI3VX1
Xg16948__7482 n_83 n_75 n_140 n_180 gnd3i! vdd3i! / ON21JI3VX1
Xg16870__5526 n_244 npg1_phase_up_count<0> n_66 n_277 gnd3i! vdd3i! / 
+ ON21JI3VX1
Xg16729__1617 n_320 npg1_freq_count<9> n_394 n_406 gnd3i! vdd3i! / ON21JI3VX1
Xg16611__9945 n_431 n_353 n_473 n_481 gnd3i! vdd3i! / ON21JI3VX1
Xg16810__6131 n_158 n_11 n_312 n_324 gnd3i! vdd3i! / ON21JI3VX1
Xg16895__7410 n_58 conf0<19> conf0<18> n_239 gnd3i! vdd3i! / ON21JI3VX1
Xg16800__6783 n_305 n_3 n_0 n_334 gnd3i! vdd3i! / ON21JI3VX1
Xg16867__6260 n_245 npg1_DOWN_count<4> n_55 n_270 gnd3i! vdd3i! / ON21JI3VX1
Xg16708__6417 n_355 n_351 n_400 n_410 gnd3i! vdd3i! / ON21JI3VX1
Xg16889__9315 n_211 n_139 n_744 n_247 gnd3i! vdd3i! / ON21JI3VX1
Xg16827__7410 n_248 n_117 n_215 n_310 gnd3i! vdd3i! / ON21JI3VX1
Xg16930__6260 n_136 n_118 n_90 n_206 gnd3i! vdd3i! / ON21JI3VX1
Xg16977__6131 n_44 conf1<10> n_86 n_154 gnd3i! vdd3i! / ON21JI3VX1
Xg16811__1881 n_279 n_254 npg1_phase_down_count<2> n_323 gnd3i! vdd3i! / 
+ ON21JI3VX1
Xg16797__4319 n_251 n_127 n_323 n_337 gnd3i! vdd3i! / ON21JI3VX1
Xspi1_Rx_count_reg[0] CTS_8 spi1_n_2088 spi1_Rx_count<0> FE_OFN30_SPI_CS 
+ gnd3i! vdd3i! / DFRRQJI3VX4
Xnpg1_phase_down_count_reg[0] CTS_4 n_301 npg1_phase_down_count<0> 
+ FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX4
Xnpg1_OFF_count_reg[9] CTS_2 n_479 npg1_OFF_count<9> FE_OFN33_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX4
Xnpg1_ON_count_reg[7] CTS_4 n_472 npg1_ON_count<7> FE_PHN271_n_32 gnd3i! 
+ vdd3i! / DFRRQJI3VX4
Xnpg1_phase_up_count_reg[2] CTS_4 n_332 npg1_phase_up_count<2> FE_PHN271_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX4
Xnpg1_phase_up_count_reg[1] CTS_4 n_314 npg1_phase_up_count<1> FE_PHN271_n_32 
+ gnd3i! vdd3i! / DFRRQJI3VX4
Xnpg1_phase_down_count_reg[2] CTS_4 n_337 npg1_phase_down_count<2> 
+ FE_PHN271_n_32 gnd3i! vdd3i! / DFRRQJI3VX4
Xg16860__6417 n_739 FE_OFN50_npg1_phase_up_state npg1_pulse_start n_281 gnd3i! 
+ vdd3i! / AO21JI3VX1
Xg16668__6417 n_403 npg1_OFF_count<0> n_432 n_441 gnd3i! vdd3i! / AO21JI3VX1
Xg16975__8246 n_25 conf0<12> n_96 n_156 gnd3i! vdd3i! / AO21JI3VX1
Xg16781__4733 npg1_freq_count<0> n_11 n_340 n_352 gnd3i! vdd3i! / AO21JI3VX1
Xg16672__6260 n_426 n_366 n_405 n_444 gnd3i! vdd3i! / AO21JI3VX1
Xg16669__5477 n_426 n_213 n_405 n_447 gnd3i! vdd3i! / AO21JI3VX1
Xg16996__4319 npg1_UP_count<1> n_26 n_119 n_131 gnd3i! vdd3i! / AO21JI3VX1
Xg17150__2398 n_70 n_78 n_100 n_8 gnd3i! vdd3i! / AO21JI3VX1
Xg11746__5122 FE_OFN10_up_switches_21 FE_OFN9_up_switches_23 
+ FE_OFN8_up_switches_24 n_642 gnd3i! vdd3i! / OR3JI3VX1
Xg11745__1705 n_638 FE_OFN26_up_switches_3 FE_OFN27_up_switches_2 n_643 gnd3i! 
+ vdd3i! / OR3JI3VX1
Xg16910__8246 n_176 n_171 n_177 n_236 gnd3i! vdd3i! / OR3JI3VX1
Xg16967__3680 n_152 n_84 n_107 n_167 gnd3i! vdd3i! / OR3JI3VX1
Xg16927__5477 n_167 n_147 n_143 n_209 gnd3i! vdd3i! / OR3JI3VX1
Xspi1_g942__7482 spi1_n_2001 spi1_n_2014 spi1_n_2015 spi1_n_1998 gnd3i! vdd3i! 
+ / NO3JI3VX0
Xg16703__2883 n_405 n_395 n_11 n_426 gnd3i! vdd3i! / NO3JI3VX0
Xg16905__3680 n_139 n_181 n_175 n_232 gnd3i! vdd3i! / NO3JI3VX0
Xg16961__5107 n_112 n_118 n_154 n_173 gnd3i! vdd3i! / NO3JI3VX0
Xg16944__6131 n_123 n_1 n_128 n_183 gnd3i! vdd3i! / NO3I1JI3VX1
Xg2__6417 n_274 n_264 n_291 n_10 gnd3i! vdd3i! / NO3I1JI3VX1
Xg16929__5107 n_4 n_124 n_168 n_207 gnd3i! vdd3i! / NO3I1JI3VX1
Xg16904__6783 n_744 n_144 n_166 n_233 gnd3i! vdd3i! / NO3I1JI3VX1
Xg16891__2883 n_215 n_221 n_209 n_252 gnd3i! vdd3i! / NO3I1JI3VX1
Xg17170 n_510 ele2<23> FE_OFN50_npg1_phase_up_state ele1<23> 
+ FE_OFN9_up_switches_23 gnd3i! vdd3i! / AO22JI3VX1
Xg16659__7482 n_430 n_194 n_423 npg1_UP_accumulator<0> n_454 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16660__4733 n_430 n_259 n_423 npg1_UP_accumulator<1> n_453 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16661__6161 n_430 n_329 n_423 npg1_UP_accumulator<2> n_452 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16662__9315 n_430 n_373 n_423 npg1_UP_accumulator<3> n_451 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16663__9945 n_430 n_420 n_423 npg1_UP_accumulator<4> n_450 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16610__9315 n_430 n_467 n_423 npg1_UP_accumulator<5> n_482 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16593__6131 n_430 n_486 n_423 npg1_UP_accumulator<6> n_490 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16588__5122 n_494 n_430 n_423 npg1_UP_accumulator<7> n_495 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16580__5526 n_498 n_430 n_423 npg1_UP_accumulator<8> n_503 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16575__6260 n_501 n_430 n_423 npg1_UP_accumulator<9> n_506 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg17169 n_510 ele2<24> FE_OFN50_npg1_phase_up_state ele1<24> 
+ FE_OFN8_up_switches_24 gnd3i! vdd3i! / AO22JI3VX1
Xg11850__5477 n_510 ele2<21> FE_OFN50_npg1_phase_up_state ele1<21> 
+ FE_OFN10_up_switches_21 gnd3i! vdd3i! / AO22JI3VX1
Xg16748__2346 n_356 n_192 n_339 FE_PHN401_npg1_DOWN_accumulator_0 n_383 gnd3i! 
+ vdd3i! / AO22JI3VX1
Xg16749__1666 n_356 n_257 n_339 npg1_DOWN_accumulator<1> n_382 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16750__7410 n_356 n_327 n_339 npg1_DOWN_accumulator<2> n_381 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16723__6260 n_356 n_375 n_339 npg1_DOWN_accumulator<3> n_402 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16681__1705 n_356 n_422 n_339 npg1_DOWN_accumulator<4> n_434 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16609__6161 n_356 n_465 n_339 npg1_DOWN_accumulator<5> n_483 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16594__1881 n_356 n_488 n_339 npg1_DOWN_accumulator<6> n_489 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16587__1705 n_492 n_356 n_339 npg1_DOWN_accumulator<7> n_496 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16579__8428 n_500 n_356 n_339 npg1_DOWN_accumulator<8> n_504 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16576__4319 n_502 n_356 n_339 npg1_DOWN_accumulator<9> n_505 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg11802__5115 n_509 ele2<1> FE_OFN57_npg1_phase_up_state ele1<1> 
+ FE_OFN28_up_switches_1 gnd3i! vdd3i! / AO22JI3VX1
Xg11847__1666 n_509 ele2<9> FE_OFN57_npg1_phase_up_state ele1<9> 
+ FE_OFN20_up_switches_9 gnd3i! vdd3i! / AO22JI3VX1
Xg11792__6783 n_509 ele2<8> FE_OFN57_npg1_phase_up_state ele1<8> 
+ FE_OFN21_up_switches_8 gnd3i! vdd3i! / AO22JI3VX1
Xg11803__7482 n_509 ele2<0> FE_OFN57_npg1_phase_up_state ele1<0> 
+ FE_OFN29_up_switches_0 gnd3i! vdd3i! / AO22JI3VX1
Xg11801__1881 n_509 ele2<2> FE_OFN57_npg1_phase_up_state ele1<2> 
+ FE_OFN27_up_switches_2 gnd3i! vdd3i! / AO22JI3VX1
Xg11800__6131 n_509 ele2<3> FE_OFN57_npg1_phase_up_state ele1<3> 
+ FE_OFN26_up_switches_3 gnd3i! vdd3i! / AO22JI3VX1
Xg11799__7098 n_509 ele2<4> FE_OFN57_npg1_phase_up_state ele1<4> 
+ FE_OFN25_up_switches_4 gnd3i! vdd3i! / AO22JI3VX1
Xg11798__8246 n_509 ele2<5> FE_OFN57_npg1_phase_up_state ele1<5> 
+ FE_OFN24_up_switches_5 gnd3i! vdd3i! / AO22JI3VX1
Xg11843__9315 n_509 ele2<10> FE_OFN57_npg1_phase_up_state ele1<10> 
+ FE_OFN19_up_switches_10 gnd3i! vdd3i! / AO22JI3VX1
Xg11844__9945 n_509 ele2<11> FE_OFN57_npg1_phase_up_state ele1<11> 
+ FE_OFN18_up_switches_11 gnd3i! vdd3i! / AO22JI3VX1
Xg11797__5122 n_509 ele2<6> FE_OFN57_npg1_phase_up_state ele1<6> 
+ FE_OFN23_up_switches_6 gnd3i! vdd3i! / AO22JI3VX1
Xg11789__4319 n_509 ele2<7> FE_OFN57_npg1_phase_up_state ele1<7> 
+ FE_OFN22_up_switches_7 gnd3i! vdd3i! / AO22JI3VX1
Xg11846__2346 n_509 ele2<12> FE_OFN57_npg1_phase_up_state ele1<12> 
+ FE_OFN17_up_switches_12 gnd3i! vdd3i! / AO22JI3VX1
Xg11848__7410 n_509 ele2<13> FE_OFN57_npg1_phase_up_state ele1<13> 
+ FE_OFN16_up_switches_13 gnd3i! vdd3i! / AO22JI3VX1
Xg11796__1705 n_510 ele2<20> FE_OFN50_npg1_phase_up_state ele1<20> 
+ FE_OFN11_up_switches_20 gnd3i! vdd3i! / AO22JI3VX1
Xg16679__1617 n_413 n_288 n_403 npg1_OFF_count<5> n_436 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16676__5526 n_413 n_346 n_403 npg1_OFF_count<6> n_439 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16677__6783 n_413 n_367 n_403 npg1_OFF_count<7> n_438 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16710__2398 n_386 n_319 n_371 npg1_freq_count<8> n_408 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16680__2802 n_426 n_360 n_405 npg1_ON_count<5> n_435 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16636__8428 n_447 npg1_ON_count<4> n_426 n_317 n_470 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16678__3680 n_426 n_187 n_405 npg1_ON_count<1> n_437 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16675__8428 n_426 n_230 n_405 npg1_ON_count<2> n_440 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16779__5115 n_319 n_246 FE_PHN407_npg1_freq_count_5 n_11 n_354 gnd3i! vdd3i! 
+ / AO22JI3VX1
Xg16762__5526 n_319 n_316 npg1_freq_count<6> n_11 n_370 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16753__2398 n_356 n_189 n_339 npg1_DOWN_count<1> n_378 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16746__9945 n_356 n_255 n_339 npg1_DOWN_count<2> n_385 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16747__2883 n_356 n_293 n_339 npg1_DOWN_count<3> n_384 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16664__2883 n_430 n_190 n_423 npg1_UP_count<1> n_449 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16657__1881 n_430 n_292 n_423 npg1_UP_count<3> n_456 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16665__2346 n_430 n_260 n_423 npg1_UP_count<2> n_448 gnd3i! vdd3i! / 
+ AO22JI3VX1
Xg16924__1666 n_141 n_84 n_143 n_93 n_212 gnd3i! vdd3i! / AO22JI3VX1
Xg16893__1666 n_183 n_202 n_217 n_199 n_250 gnd3i! vdd3i! / AN31JI3VX1
Xg16764__3680 n_64 n_120 n_334 n_63 n_368 gnd3i! vdd3i! / AN31JI3VX1
Xg16771__8246 n_73 n_238 n_310 n_91 n_358 gnd3i! vdd3i! / AN31JI3VX1
Xspi1_g988__2883 IC_addr<0> spi1_Rx_data_temp<38> spi1_n_2014 gnd3i! vdd3i! / 
+ EO2JI3VX0
Xspi1_g989__2346 IC_addr<1> spi1_Rx_data_temp<39> spi1_n_2015 gnd3i! vdd3i! / 
+ EO2JI3VX0
Xg16765__1617 n_347 npg1_OFF_count<7> n_367 gnd3i! vdd3i! / EO2JI3VX0
Xg16907__2802 n_204 npg1_ON_count<2> n_230 gnd3i! vdd3i! / EO2JI3VX0
Xg16850__5115 n_266 npg1_DOWN_count<3> n_293 gnd3i! vdd3i! / EO2JI3VX0
Xg16851__7482 n_267 npg1_UP_count<3> n_292 gnd3i! vdd3i! / EO2JI3VX0
Xg16840__6783 n_235 n_145 n_303 gnd3i! vdd3i! / EO2JI3VX0
Xg16903__5526 n_146 n_96 n_234 gnd3i! vdd3i! / EO2JI3VX0
Xg16879__5122 conf1<1> npg1_UP_accumulator<1> n_193 n_258 n_259 gnd3i! vdd3i! 
+ / FAJI3VX1
Xg16757__8428 conf1<3> npg1_UP_accumulator<3> n_328 n_372 n_373 gnd3i! vdd3i! 
+ / FAJI3VX1
Xg16807__5122 conf1<2> npg1_UP_accumulator<2> n_258 n_328 n_329 gnd3i! vdd3i! 
+ / FAJI3VX1
Xg16639__3680 conf1<5> npg1_UP_accumulator<5> n_419 n_466 n_467 gnd3i! vdd3i! 
+ / FAJI3VX1
Xg16697__4733 conf1<4> npg1_UP_accumulator<4> n_372 n_419 n_420 gnd3i! vdd3i! 
+ / FAJI3VX1
Xg16589__8246 conf1<7> npg1_UP_accumulator<7> n_485 n_493 n_494 gnd3i! vdd3i! 
+ / FAJI3VX1
Xg16596__7482 conf1<6> npg1_UP_accumulator<6> n_466 n_485 n_486 gnd3i! vdd3i! 
+ / FAJI3VX1
Xg16584__2802 conf1<8> npg1_UP_accumulator<8> n_493 n_497 n_498 gnd3i! vdd3i! 
+ / FAJI3VX1
Xg16880__8246 conf1<1> npg1_DOWN_accumulator<1> n_191 n_256 n_257 gnd3i! 
+ vdd3i! / FAJI3VX1
Xg16756__4319 conf1<3> npg1_DOWN_accumulator<3> n_326 n_374 n_375 gnd3i! 
+ vdd3i! / FAJI3VX1
Xg16808__8246 conf1<2> npg1_DOWN_accumulator<2> n_256 n_326 n_327 gnd3i! 
+ vdd3i! / FAJI3VX1
Xg16640__1617 conf1<5> npg1_DOWN_accumulator<5> n_421 n_464 n_465 gnd3i! 
+ vdd3i! / FAJI3VX1
Xg16696__7482 conf1<4> npg1_DOWN_accumulator<4> n_374 n_421 n_422 gnd3i! 
+ vdd3i! / FAJI3VX1
Xg16590__7098 conf1<7> npg1_DOWN_accumulator<7> n_487 n_491 n_492 gnd3i! 
+ vdd3i! / FAJI3VX1
Xg16595__5115 conf1<6> npg1_DOWN_accumulator<6> n_464 n_487 n_488 gnd3i! 
+ vdd3i! / FAJI3VX1
Xg16583__1617 conf1<8> npg1_DOWN_accumulator<8> n_491 n_499 n_500 gnd3i! 
+ vdd3i! / FAJI3VX1
Xg16698__6161 n_31 npg1_DOWN_accumulator<8> n_376 n_417 n_418 gnd3i! vdd3i! / 
+ FAJI3VX1
Xg16755__6260 n_30 npg1_DOWN_accumulator<7> n_290 n_376 n_377 gnd3i! vdd3i! / 
+ FAJI3VX1
XFE_PHC410_spi1_n_1763 spi1_n_1763 FE_PHN410_spi1_n_1763 gnd3i! vdd3i! / 
+ BUJI3VX0
XFE_PHC404_spi1_Rx_count_4 spi1_Rx_count<4> FE_PHN404_spi1_Rx_count_4 gnd3i! 
+ vdd3i! / BUJI3VX0
XFE_PHC416_SPI_MOSI SPI_MOSI FE_PHN416_SPI_MOSI gnd3i! vdd3i! / BUJI3VX0
XFE_PHC448_n_32 FE_PHN428_n_32 FE_PHN448_n_32 gnd3i! vdd3i! / BUJI3VX0
XFE_PHC429_n_32 FE_PHN427_n_32 FE_PHN429_n_32 gnd3i! vdd3i! / BUJI3VX0
XFE_PHC423_n_32 FE_PHN424_n_32 FE_PHN423_n_32 gnd3i! vdd3i! / BUJI3VX0
XFE_PHC424_n_32 FE_PHN425_n_32 FE_PHN424_n_32 gnd3i! vdd3i! / BUJI3VX0
XFE_PHC425_n_32 FE_PHN426_n_32 FE_PHN425_n_32 gnd3i! vdd3i! / BUJI3VX0
XFE_PHC426_n_32 n_32 FE_PHN426_n_32 gnd3i! vdd3i! / BUJI3VX0
XFE_PHC419_porborn FE_PHN420_porborn FE_PHN419_porborn gnd3i! vdd3i! / BUJI3VX0
XFE_PHC420_porborn FE_PHN417_porborn FE_PHN420_porborn gnd3i! vdd3i! / BUJI3VX0
XFE_PHC417_porborn FE_PHN408_porborn FE_PHN417_porborn gnd3i! vdd3i! / BUJI3VX0
XFE_PHC408_porborn porborn FE_PHN408_porborn gnd3i! vdd3i! / BUJI3VX0
XFE_PHC406_spi1_Rx_count_1 spi1_Rx_count<1> FE_PHN406_spi1_Rx_count_1 gnd3i! 
+ vdd3i! / BUJI3VX0
XFE_PHC412_spi1_Rx_data_temp_36 spi1_Rx_data_temp<36> 
+ FE_PHN412_spi1_Rx_data_temp_36 gnd3i! vdd3i! / BUJI3VX0
XFE_PHC414_spi1_Rx_data_temp_35 spi1_Rx_data_temp<35> 
+ FE_PHN414_spi1_Rx_data_temp_35 gnd3i! vdd3i! / BUJI3VX0
XFE_PHC401_npg1_DOWN_accumulator_0 npg1_DOWN_accumulator<0> 
+ FE_PHN401_npg1_DOWN_accumulator_0 gnd3i! vdd3i! / BUJI3VX0
XFE_PHC405_npg1_OFF_count_0 npg1_OFF_count<0> FE_PHN405_npg1_OFF_count_0 
+ gnd3i! vdd3i! / BUJI3VX0
XFE_PHC397_npg1_OFF_count_3 npg1_OFF_count<3> FE_PHN397_npg1_OFF_count_3 
+ gnd3i! vdd3i! / BUJI3VX0
XFE_PHC403_conf0_13 conf0<13> FE_PHN403_conf0_13 gnd3i! vdd3i! / BUJI3VX0
XFE_PHC402_conf0_12 conf0<12> FE_PHN402_conf0_12 gnd3i! vdd3i! / BUJI3VX0
XFE_PHC400_conf0_14 conf0<14> FE_PHN400_conf0_14 gnd3i! vdd3i! / BUJI3VX0
XFE_PHC398_npg1_freq_count_3 npg1_freq_count<3> FE_PHN398_npg1_freq_count_3 
+ gnd3i! vdd3i! / BUJI3VX0
XFE_PHC407_npg1_freq_count_5 npg1_freq_count<5> FE_PHN407_npg1_freq_count_5 
+ gnd3i! vdd3i! / BUJI3VX0
XFE_PHC399_npg1_freq_count_10 npg1_freq_count<10> FE_PHN399_npg1_freq_count_10 
+ gnd3i! vdd3i! / BUJI3VX0
XFE_PHC409_n_442 n_442 FE_PHN409_n_442 gnd3i! vdd3i! / BUJI3VX0
XFE_PHC411_n_391 n_391 FE_PHN411_n_391 gnd3i! vdd3i! / BUJI3VX0
Xg16682__5122 n_417 npg1_DOWN_accumulator<9> conf0<17> n_433 gnd3i! vdd3i! / 
+ EN3JI3VX1
Xg17013__9315 npg1_on_off_ctrl<1> npg1_on_off_ctrl<2> npg1_on_off_ctrl<0> 
+ n_134 gnd3i! vdd3i! / NO3I2JI3VX1
Xg16787__1666 n_338 FE_OFN52_enable n_321 n_356 gnd3i! vdd3i! / NO3I2JI3VX1
Xspi1_g930__1705 spi1_n_1929 FE_PHN404_spi1_Rx_count_4 spi1_n_1926 spi1_n_1924 
+ gnd3i! vdd3i! / OA21JI3VX1
Xg16925__7410 n_137 n_106 n_103 n_211 gnd3i! vdd3i! / OA21JI3VX1
Xg16936__6783 npg1_UP_accumulator<0> conf1<0> n_193 n_194 gnd3i! vdd3i! / 
+ HAJI3VX1
Xspi1_g933__8246 spi1_n_2000 spi1_Rx_count<3> spi1_n_1929 spi1_n_1962 gnd3i! 
+ vdd3i! / HAJI3VX1
Xspi1_g943__4733 spi1_n_2018 spi1_Rx_count<2> spi1_n_2000 spi1_n_1999 gnd3i! 
+ vdd3i! / HAJI3VX1
Xg16937__3680 npg1_DOWN_accumulator<0> conf1<0> n_191 n_192 gnd3i! vdd3i! / 
+ HAJI3VX1
Xg16788__7410 n_287 npg1_OFF_count<6> n_347 n_346 gnd3i! vdd3i! / HAJI3VX1
Xg16854__9315 n_216 npg1_OFF_count<5> n_287 n_288 gnd3i! vdd3i! / HAJI3VX1
Xg16769__1705 n_304 npg1_ON_count<5> n_365 n_360 gnd3i! vdd3i! / HAJI3VX1
Xg16940__1705 npg1_ON_count<1> npg1_ON_count<0> n_204 n_187 gnd3i! vdd3i! / 
+ HAJI3VX1
Xg16939__2802 npg1_DOWN_count<1> npg1_DOWN_count<0> n_188 n_189 gnd3i! vdd3i! 
+ / HAJI3VX1
Xg16881__7098 n_188 npg1_DOWN_count<2> n_266 n_255 gnd3i! vdd3i! / HAJI3VX1
Xg16938__1617 npg1_UP_count<1> npg1_UP_count<0> n_205 n_190 gnd3i! vdd3i! / 
+ HAJI3VX1
Xg16878__1705 n_205 npg1_UP_count<2> n_267 n_260 gnd3i! vdd3i! / HAJI3VX1
XFE_PHC275_SPI_CS SPI_CS FE_PHN275_SPI_CS gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC348_spi1_conf1_meta_1 spi1_conf1_meta<1> FE_PHN348_spi1_conf1_meta_1 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC293_spi1_conf1_meta_3 spi1_conf1_meta<3> FE_PHN293_spi1_conf1_meta_3 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC303_spi1_conf1_meta_6 spi1_conf1_meta<6> FE_PHN303_spi1_conf1_meta_6 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC296_spi1_ele2_meta_31 spi1_ele2_meta<31> FE_PHN296_spi1_ele2_meta_31 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC338_spi1_ele2_meta_30 spi1_ele2_meta<30> FE_PHN338_spi1_ele2_meta_30 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC276_spi1_ele2_meta_29 spi1_ele2_meta<29> FE_PHN276_spi1_ele2_meta_29 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC333_spi1_ele2_meta_28 spi1_ele2_meta<28> FE_PHN333_spi1_ele2_meta_28 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC340_spi1_ele2_meta_27 spi1_ele2_meta<27> FE_PHN340_spi1_ele2_meta_27 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC366_spi1_conf0_meta_20 spi1_conf0_meta<20> FE_PHN366_spi1_conf0_meta_20 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC346_spi1_conf0_meta_19 spi1_conf0_meta<19> FE_PHN346_spi1_conf0_meta_19 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC396_spi1_conf1_meta_5 spi1_conf1_meta<5> FE_PHN396_spi1_conf1_meta_5 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC395_spi1_ele2_meta_8 spi1_ele2_meta<8> FE_PHN395_spi1_ele2_meta_8 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC394_spi1_conf1_meta_9 spi1_conf1_meta<9> FE_PHN394_spi1_conf1_meta_9 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC393_spi1_ele2_meta_6 spi1_ele2_meta<6> FE_PHN393_spi1_ele2_meta_6 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC392_spi1_ele1_meta_8 spi1_ele1_meta<8> FE_PHN392_spi1_ele1_meta_8 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC391_spi1_ele1_meta_19 spi1_ele1_meta<19> FE_PHN391_spi1_ele1_meta_19 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC390_spi1_conf0_meta_21 spi1_conf0_meta<21> FE_PHN390_spi1_conf0_meta_21 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC389_spi1_conf1_meta_7 spi1_conf1_meta<7> FE_PHN389_spi1_conf1_meta_7 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC388_spi1_ele2_meta_26 spi1_ele2_meta<26> FE_PHN388_spi1_ele2_meta_26 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC387_spi1_conf1_meta_4 spi1_conf1_meta<4> FE_PHN387_spi1_conf1_meta_4 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC386_spi1_conf0_meta_0 spi1_conf0_meta<0> FE_PHN386_spi1_conf0_meta_0 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC385_spi1_ele2_meta_14 spi1_ele2_meta<14> FE_PHN385_spi1_ele2_meta_14 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC384_spi1_conf1_meta_16 spi1_conf1_meta<16> FE_PHN384_spi1_conf1_meta_16 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC383_spi1_ele2_meta_22 spi1_ele2_meta<22> FE_PHN383_spi1_ele2_meta_22 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC382_spi1_ele1_meta_2 spi1_ele1_meta<2> FE_PHN382_spi1_ele1_meta_2 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC381_spi1_ele1_meta_24 spi1_ele1_meta<24> FE_PHN381_spi1_ele1_meta_24 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC380_spi1_ele2_meta_10 spi1_ele2_meta<10> FE_PHN380_spi1_ele2_meta_10 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC379_spi1_conf0_meta_30 spi1_conf0_meta<30> FE_PHN379_spi1_conf0_meta_30 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC378_spi1_conf1_meta_17 spi1_conf1_meta<17> FE_PHN378_spi1_conf1_meta_17 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC377_spi1_conf0_meta_18 spi1_conf0_meta<18> FE_PHN377_spi1_conf0_meta_18 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC376_spi1_conf1_meta_2 spi1_conf1_meta<2> FE_PHN376_spi1_conf1_meta_2 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC375_spi1_ele1_meta_31 spi1_ele1_meta<31> FE_PHN375_spi1_ele1_meta_31 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC374_spi1_conf1_meta_10 spi1_conf1_meta<10> FE_PHN374_spi1_conf1_meta_10 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC373_spi1_conf0_meta_27 spi1_conf0_meta<27> FE_PHN373_spi1_conf0_meta_27 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC372_spi1_conf1_meta_12 spi1_conf1_meta<12> FE_PHN372_spi1_conf1_meta_12 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC371_spi1_ele1_meta_29 spi1_ele1_meta<29> FE_PHN371_spi1_ele1_meta_29 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC370_spi1_ele1_meta_16 spi1_ele1_meta<16> FE_PHN370_spi1_ele1_meta_16 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC369_spi1_conf0_meta_5 spi1_conf0_meta<5> FE_PHN369_spi1_conf0_meta_5 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC368_spi1_ele2_meta_16 spi1_ele2_meta<16> FE_PHN368_spi1_ele2_meta_16 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC367_spi1_conf0_meta_8 spi1_conf0_meta<8> FE_PHN367_spi1_conf0_meta_8 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC365_spi1_conf0_meta_13 spi1_conf0_meta<13> FE_PHN365_spi1_conf0_meta_13 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC364_spi1_conf0_meta_24 spi1_conf0_meta<24> FE_PHN364_spi1_conf0_meta_24 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC363_spi1_ele1_meta_22 spi1_ele1_meta<22> FE_PHN363_spi1_ele1_meta_22 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC362_spi1_ele1_meta_28 spi1_ele1_meta<28> FE_PHN362_spi1_ele1_meta_28 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC361_spi1_conf1_meta_11 spi1_conf1_meta<11> FE_PHN361_spi1_conf1_meta_11 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC360_spi1_conf0_meta_14 spi1_conf0_meta<14> FE_PHN360_spi1_conf0_meta_14 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC359_spi1_ele1_meta_23 spi1_ele1_meta<23> FE_PHN359_spi1_ele1_meta_23 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC358_spi1_ele2_meta_7 spi1_ele2_meta<7> FE_PHN358_spi1_ele2_meta_7 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC357_spi1_conf0_meta_9 spi1_conf0_meta<9> FE_PHN357_spi1_conf0_meta_9 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC356_spi1_conf1_meta_21 spi1_conf1_meta<21> FE_PHN356_spi1_conf1_meta_21 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC355_spi1_conf1_meta_23 spi1_conf1_meta<23> FE_PHN355_spi1_conf1_meta_23 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC354_spi1_ele1_meta_17 spi1_ele1_meta<17> FE_PHN354_spi1_ele1_meta_17 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC353_spi1_conf0_meta_7 spi1_conf0_meta<7> FE_PHN353_spi1_conf0_meta_7 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC352_spi1_conf1_meta_22 spi1_conf1_meta<22> FE_PHN352_spi1_conf1_meta_22 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC351_spi1_conf1_meta_13 spi1_conf1_meta<13> FE_PHN351_spi1_conf1_meta_13 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC350_spi1_ele1_meta_6 spi1_ele1_meta<6> FE_PHN350_spi1_ele1_meta_6 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC349_spi1_ele1_meta_0 spi1_ele1_meta<0> FE_PHN349_spi1_ele1_meta_0 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC347_spi1_conf0_meta_26 spi1_conf0_meta<26> FE_PHN347_spi1_conf0_meta_26 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC298_spi1_conf0_meta_22 spi1_conf0_meta<22> FE_PHN298_spi1_conf0_meta_22 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC345_spi1_conf0_meta_28 spi1_conf0_meta<28> FE_PHN345_spi1_conf0_meta_28 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC344_spi1_ele1_meta_26 spi1_ele1_meta<26> FE_PHN344_spi1_ele1_meta_26 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC343_spi1_ele2_meta_3 spi1_ele2_meta<3> FE_PHN343_spi1_ele2_meta_3 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC342_spi1_conf0_meta_25 spi1_conf0_meta<25> FE_PHN342_spi1_conf0_meta_25 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC341_spi1_ele2_meta_15 spi1_ele2_meta<15> FE_PHN341_spi1_ele2_meta_15 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC337_spi1_ele1_meta_7 spi1_ele1_meta<7> FE_PHN337_spi1_ele1_meta_7 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC336_spi1_ele2_meta_24 spi1_ele2_meta<24> FE_PHN336_spi1_ele2_meta_24 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC335_spi1_ele1_meta_30 spi1_ele1_meta<30> FE_PHN335_spi1_ele1_meta_30 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC334_spi1_conf0_meta_6 spi1_conf0_meta<6> FE_PHN334_spi1_conf0_meta_6 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC332_spi1_ele1_meta_5 spi1_ele1_meta<5> FE_PHN332_spi1_ele1_meta_5 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC331_spi1_ele2_meta_12 spi1_ele2_meta<12> FE_PHN331_spi1_ele2_meta_12 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC330_spi1_ele1_meta_1 spi1_ele1_meta<1> FE_PHN330_spi1_ele1_meta_1 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC328_spi1_ele1_meta_20 spi1_ele1_meta<20> FE_PHN328_spi1_ele1_meta_20 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC327_spi1_ele1_meta_25 spi1_ele1_meta<25> FE_PHN327_spi1_ele1_meta_25 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC326_spi1_ele1_meta_4 spi1_ele1_meta<4> FE_PHN326_spi1_ele1_meta_4 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC325_spi1_ele2_meta_11 spi1_ele2_meta<11> FE_PHN325_spi1_ele2_meta_11 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC324_spi1_ele2_meta_2 spi1_ele2_meta<2> FE_PHN324_spi1_ele2_meta_2 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC323_spi1_ele1_meta_13 spi1_ele1_meta<13> FE_PHN323_spi1_ele1_meta_13 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC322_spi1_ele1_meta_3 spi1_ele1_meta<3> FE_PHN322_spi1_ele1_meta_3 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC321_spi1_ele1_meta_18 spi1_ele1_meta<18> FE_PHN321_spi1_ele1_meta_18 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC320_spi1_ele2_meta_5 spi1_ele2_meta<5> FE_PHN320_spi1_ele2_meta_5 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC319_spi1_ele2_meta_23 spi1_ele2_meta<23> FE_PHN319_spi1_ele2_meta_23 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC318_spi1_conf0_meta_29 spi1_conf0_meta<29> FE_PHN318_spi1_conf0_meta_29 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC317_spi1_conf0_meta_12 spi1_conf0_meta<12> FE_PHN317_spi1_conf0_meta_12 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC316_spi1_ele1_meta_21 spi1_ele1_meta<21> FE_PHN316_spi1_ele1_meta_21 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC315_spi1_ele2_meta_20 spi1_ele2_meta<20> FE_PHN315_spi1_ele2_meta_20 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC313_spi1_ele2_meta_25 spi1_ele2_meta<25> FE_PHN313_spi1_ele2_meta_25 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC312_spi1_ele2_meta_13 spi1_ele2_meta<13> FE_PHN312_spi1_ele2_meta_13 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC311_spi1_ele2_meta_21 spi1_ele2_meta<21> FE_PHN311_spi1_ele2_meta_21 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC310_spi1_conf0_meta_10 spi1_conf0_meta<10> FE_PHN310_spi1_conf0_meta_10 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC309_spi1_ele1_meta_27 spi1_ele1_meta<27> FE_PHN309_spi1_ele1_meta_27 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC308_spi1_ele1_meta_9 spi1_ele1_meta<9> FE_PHN308_spi1_ele1_meta_9 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC307_spi1_conf0_meta_17 spi1_conf0_meta<17> FE_PHN307_spi1_conf0_meta_17 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC306_spi1_ele2_meta_19 spi1_ele2_meta<19> FE_PHN306_spi1_ele2_meta_19 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC305_spi1_conf0_meta_1 spi1_conf0_meta<1> FE_PHN305_spi1_conf0_meta_1 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC304_spi1_conf0_meta_16 spi1_conf0_meta<16> FE_PHN304_spi1_conf0_meta_16 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC302_spi1_conf0_meta_23 spi1_conf0_meta<23> FE_PHN302_spi1_conf0_meta_23 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC301_spi1_ele1_meta_15 spi1_ele1_meta<15> FE_PHN301_spi1_ele1_meta_15 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC300_spi1_ele2_meta_9 spi1_ele2_meta<9> FE_PHN300_spi1_ele2_meta_9 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC299_spi1_ele2_meta_1 spi1_ele2_meta<1> FE_PHN299_spi1_ele2_meta_1 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC297_spi1_ele1_meta_10 spi1_ele1_meta<10> FE_PHN297_spi1_ele1_meta_10 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC295_spi1_ele2_meta_18 spi1_ele2_meta<18> FE_PHN295_spi1_ele2_meta_18 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC290_spi1_ele2_meta_0 spi1_ele2_meta<0> FE_PHN290_spi1_ele2_meta_0 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC289_spi1_ele2_meta_4 spi1_ele2_meta<4> FE_PHN289_spi1_ele2_meta_4 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC288_spi1_conf0_meta_31 spi1_conf0_meta<31> FE_PHN288_spi1_conf0_meta_31 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC286_spi1_conf0_meta_15 spi1_conf0_meta<15> FE_PHN286_spi1_conf0_meta_15 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC285_spi1_ele1_meta_14 spi1_ele1_meta<14> FE_PHN285_spi1_ele1_meta_14 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC284_spi1_conf0_meta_3 spi1_conf0_meta<3> FE_PHN284_spi1_conf0_meta_3 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC283_spi1_conf0_meta_2 spi1_conf0_meta<2> FE_PHN283_spi1_conf0_meta_2 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC281_spi1_conf0_meta_4 spi1_conf0_meta<4> FE_PHN281_spi1_conf0_meta_4 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC280_spi1_conf0_meta_11 spi1_conf0_meta<11> FE_PHN280_spi1_conf0_meta_11 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC279_spi1_ele2_meta_17 spi1_ele2_meta<17> FE_PHN279_spi1_ele2_meta_17 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC278_spi1_ele1_meta_12 spi1_ele1_meta<12> FE_PHN278_spi1_ele1_meta_12 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC277_spi1_ele1_meta_11 spi1_ele1_meta<11> FE_PHN277_spi1_ele1_meta_11 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC329_spi1_conf1_meta_8 spi1_conf1_meta<8> FE_PHN329_spi1_conf1_meta_8 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC292_spi1_conf1_meta_0 spi1_conf1_meta<0> FE_PHN292_spi1_conf1_meta_0 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC339_spi1_conf1_meta_18 spi1_conf1_meta<18> FE_PHN339_spi1_conf1_meta_18 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC294_spi1_conf1_meta_19 spi1_conf1_meta<19> FE_PHN294_spi1_conf1_meta_19 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC314_spi1_conf1_meta_15 spi1_conf1_meta<15> FE_PHN314_spi1_conf1_meta_15 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC291_npg1_pulse_aux npg1_pulse_aux FE_PHN291_npg1_pulse_aux gnd3i! 
+ vdd3i! / DLY1JI3VX1
XFE_PHC287_spi1_conf1_meta_20 spi1_conf1_meta<20> FE_PHN287_spi1_conf1_meta_20 
+ gnd3i! vdd3i! / DLY1JI3VX1
XFE_PHC282_spi1_conf1_meta_14 spi1_conf1_meta<14> FE_PHN282_spi1_conf1_meta_14 
+ gnd3i! vdd3i! / DLY1JI3VX1
Xspi1_g965__6161 spi1_n_2010 spi1_Rx_count<4> spi1_Rx_count<5> spi1_n_2001 
+ gnd3i! vdd3i! / NA3I2JI3VX1
Xg16945__1881 n_142 n_110 n_2 n_182 gnd3i! vdd3i! / NA3I2JI3VX1
Xg16872__3680 n_252 n_11 n_134 n_274 gnd3i! vdd3i! / NA3I2JI3VX1
Xg16963__4319 n_109 n_102 n_125 n_171 gnd3i! vdd3i! / NA3I2JI3VX1
Xg16916__5115 npg1_ON_count<1> npg1_ON_count<0> conf0<25> n_219 gnd3i! vdd3i! 
+ / NO22JI3VX1
Xg16978__1881 conf1<21> n_37 n_83 n_153 gnd3i! vdd3i! / NO22JI3VX1
Xspi1_g808__2802 spi1_Rx_count<5> spi1_n_1926 spi1_n_1763 gnd3i! vdd3i! / 
+ EN2JI3VX0
Xg16890__9945 npg1_freq_count<5> n_222 n_246 gnd3i! vdd3i! / EN2JI3VX0
Xg16820__6161 npg1_freq_count<6> n_241 n_316 gnd3i! vdd3i! / EN2JI3VX0
Xspi1_ele2_asyn_reg[31] SPI_CS spi1_Rx_data_temp<31> spi1_ele2_asyn<31> 
+ FE_PHN271_n_32 spi1_ele2_asyn<31> spi1_n_2271 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[30] SPI_CS spi1_Rx_data_temp<30> spi1_ele2_asyn<30> 
+ FE_PHN271_n_32 spi1_ele2_asyn<30> spi1_n_2271 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[29] SPI_CS spi1_Rx_data_temp<29> spi1_ele2_asyn<29> 
+ FE_PHN271_n_32 spi1_ele2_asyn<29> spi1_n_2271 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[28] SPI_CS spi1_Rx_data_temp<28> spi1_ele2_asyn<28> 
+ FE_PHN271_n_32 spi1_ele2_asyn<28> spi1_n_2271 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[27] SPI_CS spi1_Rx_data_temp<27> spi1_ele2_asyn<27> 
+ FE_PHN271_n_32 spi1_ele2_asyn<27> spi1_n_2271 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[26] SPI_CS spi1_Rx_data_temp<26> spi1_ele2_asyn<26> 
+ FE_PHN271_n_32 spi1_ele2_asyn<26> spi1_n_2271 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[25] SPI_CS spi1_Rx_data_temp<25> spi1_ele2_asyn<25> 
+ FE_PHN431_n_32 spi1_ele2_asyn<25> spi1_n_2271 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[24] SPI_CS spi1_Rx_data_temp<24> spi1_ele2_asyn<24> 
+ FE_PHN431_n_32 spi1_ele2_asyn<24> spi1_n_2271 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[23] SPI_CS spi1_Rx_data_temp<23> spi1_ele2_asyn<23> 
+ FE_PHN431_n_32 spi1_ele2_asyn<23> spi1_n_2271 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[22] FE_PHN254_SPI_CS spi1_Rx_data_temp<22> 
+ spi1_ele2_asyn<22> FE_OFN35_n_32 spi1_ele2_asyn<22> spi1_n_2271 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[21] FE_PHN254_SPI_CS spi1_Rx_data_temp<21> 
+ spi1_ele2_asyn<21> FE_OFN35_n_32 spi1_ele2_asyn<21> spi1_n_2271 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[20] FE_PHN254_SPI_CS spi1_Rx_data_temp<20> 
+ spi1_ele2_asyn<20> FE_OFN35_n_32 spi1_ele2_asyn<20> spi1_n_2271 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[19] FE_PHN254_SPI_CS spi1_Rx_data_temp<19> 
+ spi1_ele2_asyn<19> FE_OFN35_n_32 spi1_ele2_asyn<19> spi1_n_2271 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[18] FE_PHN254_SPI_CS spi1_Rx_data_temp<18> 
+ spi1_ele2_asyn<18> FE_OFN35_n_32 spi1_ele2_asyn<18> spi1_n_2271 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[17] FE_PHN254_SPI_CS spi1_Rx_data_temp<17> 
+ spi1_ele2_asyn<17> FE_OFN35_n_32 spi1_ele2_asyn<17> spi1_n_2271 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[16] FE_PHN254_SPI_CS spi1_Rx_data_temp<16> 
+ spi1_ele2_asyn<16> FE_OFN35_n_32 spi1_ele2_asyn<16> spi1_n_2271 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[15] FE_PHN254_SPI_CS spi1_Rx_data_temp<15> 
+ spi1_ele2_asyn<15> FE_PHN421_n_32 spi1_ele2_asyn<15> spi1_n_2271 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[14] FE_PHN254_SPI_CS spi1_Rx_data_temp<14> 
+ spi1_ele2_asyn<14> FE_PHN421_n_32 spi1_ele2_asyn<14> spi1_n_2271 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[13] FE_PHN253_SPI_CS spi1_Rx_data_temp<13> 
+ spi1_ele2_asyn<13> FE_PHN421_n_32 spi1_ele2_asyn<13> spi1_n_2271 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[12] FE_PHN253_SPI_CS spi1_Rx_data_temp<12> 
+ spi1_ele2_asyn<12> FE_PHN272_FE_OFN33_n_32 spi1_ele2_asyn<12> spi1_n_2271 
+ gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[11] FE_PHN253_SPI_CS spi1_Rx_data_temp<11> 
+ spi1_ele2_asyn<11> FE_PHN272_FE_OFN33_n_32 spi1_ele2_asyn<11> spi1_n_2271 
+ gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[10] FE_PHN253_SPI_CS spi1_Rx_data_temp<10> 
+ spi1_ele2_asyn<10> FE_PHN272_FE_OFN33_n_32 spi1_ele2_asyn<10> spi1_n_2271 
+ gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[9] FE_PHN253_SPI_CS spi1_Rx_data_temp<9> spi1_ele2_asyn<9> 
+ FE_PHN272_FE_OFN33_n_32 spi1_ele2_asyn<9> spi1_n_2271 gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[8] FE_PHN253_SPI_CS spi1_Rx_data_temp<8> spi1_ele2_asyn<8> 
+ FE_PHN272_FE_OFN33_n_32 spi1_ele2_asyn<8> spi1_n_2271 gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[7] FE_PHN253_SPI_CS spi1_Rx_data_temp<7> spi1_ele2_asyn<7> 
+ FE_PHN272_FE_OFN33_n_32 spi1_ele2_asyn<7> spi1_n_2271 gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[6] FE_PHN253_SPI_CS spi1_Rx_data_temp<6> spi1_ele2_asyn<6> 
+ FE_OFN443_FE_PHN271_n_32 spi1_ele2_asyn<6> spi1_n_2271 gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[5] FE_PHN253_SPI_CS spi1_Rx_data_temp<5> spi1_ele2_asyn<5> 
+ FE_OFN443_FE_PHN271_n_32 spi1_ele2_asyn<5> spi1_n_2271 gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[4] FE_PHN253_SPI_CS spi1_Rx_data_temp<4> spi1_ele2_asyn<4> 
+ FE_OFN443_FE_PHN271_n_32 spi1_ele2_asyn<4> spi1_n_2271 gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[3] FE_PHN253_SPI_CS spi1_Rx_data_temp<3> spi1_ele2_asyn<3> 
+ FE_PHN263_n_32 spi1_ele2_asyn<3> spi1_n_2271 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[2] FE_PHN253_SPI_CS spi1_Rx_data_temp<2> spi1_ele2_asyn<2> 
+ FE_PHN263_n_32 spi1_ele2_asyn<2> spi1_n_2271 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[1] FE_PHN253_SPI_CS spi1_Rx_data_temp<1> spi1_ele2_asyn<1> 
+ FE_PHN263_n_32 spi1_ele2_asyn<1> spi1_n_2271 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele2_asyn_reg[0] FE_PHN253_SPI_CS spi1_Rx_data_temp<0> spi1_ele2_asyn<0> 
+ FE_PHN272_FE_OFN33_n_32 spi1_ele2_asyn<0> spi1_n_2271 gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[31] SPI_CS spi1_Rx_data_temp<31> spi1_ele1_asyn<31> 
+ FE_PHN271_n_32 spi1_ele1_asyn<31> spi1_n_1930 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[30] SPI_CS spi1_Rx_data_temp<30> spi1_ele1_asyn<30> 
+ FE_PHN271_n_32 spi1_ele1_asyn<30> spi1_n_1930 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[29] SPI_CS spi1_Rx_data_temp<29> spi1_ele1_asyn<29> 
+ FE_PHN271_n_32 spi1_ele1_asyn<29> spi1_n_1930 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[28] SPI_CS spi1_Rx_data_temp<28> spi1_ele1_asyn<28> 
+ FE_PHN271_n_32 spi1_ele1_asyn<28> spi1_n_1930 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[27] SPI_CS spi1_Rx_data_temp<27> spi1_ele1_asyn<27> 
+ FE_PHN271_n_32 spi1_ele1_asyn<27> spi1_n_1930 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[26] SPI_CS spi1_Rx_data_temp<26> spi1_ele1_asyn<26> 
+ FE_PHN271_n_32 spi1_ele1_asyn<26> spi1_n_1930 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[25] SPI_CS spi1_Rx_data_temp<25> spi1_ele1_asyn<25> 
+ FE_PHN431_n_32 spi1_ele1_asyn<25> spi1_n_1930 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[24] SPI_CS spi1_Rx_data_temp<24> spi1_ele1_asyn<24> 
+ FE_PHN431_n_32 spi1_ele1_asyn<24> spi1_n_1930 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[23] SPI_CS spi1_Rx_data_temp<23> spi1_ele1_asyn<23> 
+ FE_PHN431_n_32 spi1_ele1_asyn<23> spi1_n_1930 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[22] FE_PHN254_SPI_CS spi1_Rx_data_temp<22> 
+ spi1_ele1_asyn<22> FE_OFN35_n_32 spi1_ele1_asyn<22> spi1_n_1930 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[21] FE_PHN254_SPI_CS spi1_Rx_data_temp<21> 
+ spi1_ele1_asyn<21> FE_OFN35_n_32 spi1_ele1_asyn<21> spi1_n_1930 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[20] FE_PHN254_SPI_CS spi1_Rx_data_temp<20> 
+ spi1_ele1_asyn<20> FE_OFN35_n_32 spi1_ele1_asyn<20> spi1_n_1930 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[19] SPI_CS spi1_Rx_data_temp<19> spi1_ele1_asyn<19> 
+ FE_OFN35_n_32 spi1_ele1_asyn<19> spi1_n_1930 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[18] FE_PHN254_SPI_CS spi1_Rx_data_temp<18> 
+ spi1_ele1_asyn<18> FE_OFN35_n_32 spi1_ele1_asyn<18> spi1_n_1930 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[17] FE_PHN254_SPI_CS spi1_Rx_data_temp<17> 
+ spi1_ele1_asyn<17> FE_OFN35_n_32 spi1_ele1_asyn<17> spi1_n_1930 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[16] FE_PHN254_SPI_CS spi1_Rx_data_temp<16> 
+ spi1_ele1_asyn<16> FE_OFN35_n_32 spi1_ele1_asyn<16> spi1_n_1930 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[15] FE_PHN254_SPI_CS spi1_Rx_data_temp<15> 
+ spi1_ele1_asyn<15> FE_OFN35_n_32 spi1_ele1_asyn<15> spi1_n_1930 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[14] FE_PHN253_SPI_CS spi1_Rx_data_temp<14> 
+ spi1_ele1_asyn<14> FE_PHN421_n_32 spi1_ele1_asyn<14> spi1_n_1930 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[13] FE_PHN254_SPI_CS spi1_Rx_data_temp<13> 
+ spi1_ele1_asyn<13> FE_PHN421_n_32 spi1_ele1_asyn<13> spi1_n_1930 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[12] FE_PHN253_SPI_CS spi1_Rx_data_temp<12> 
+ spi1_ele1_asyn<12> FE_PHN272_FE_OFN33_n_32 spi1_ele1_asyn<12> spi1_n_1930 
+ gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[11] FE_PHN253_SPI_CS spi1_Rx_data_temp<11> 
+ spi1_ele1_asyn<11> FE_PHN272_FE_OFN33_n_32 spi1_ele1_asyn<11> spi1_n_1930 
+ gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[10] FE_PHN253_SPI_CS spi1_Rx_data_temp<10> 
+ spi1_ele1_asyn<10> FE_PHN272_FE_OFN33_n_32 spi1_ele1_asyn<10> spi1_n_1930 
+ gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[9] FE_PHN253_SPI_CS spi1_Rx_data_temp<9> spi1_ele1_asyn<9> 
+ FE_PHN272_FE_OFN33_n_32 spi1_ele1_asyn<9> spi1_n_1930 gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[8] FE_PHN253_SPI_CS spi1_Rx_data_temp<8> spi1_ele1_asyn<8> 
+ FE_PHN272_FE_OFN33_n_32 spi1_ele1_asyn<8> spi1_n_1930 gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[7] FE_PHN253_SPI_CS spi1_Rx_data_temp<7> spi1_ele1_asyn<7> 
+ FE_OFN443_FE_PHN271_n_32 spi1_ele1_asyn<7> spi1_n_1930 gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[6] FE_PHN253_SPI_CS spi1_Rx_data_temp<6> spi1_ele1_asyn<6> 
+ FE_OFN443_FE_PHN271_n_32 spi1_ele1_asyn<6> spi1_n_1930 gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[5] FE_PHN253_SPI_CS spi1_Rx_data_temp<5> spi1_ele1_asyn<5> 
+ FE_OFN443_FE_PHN271_n_32 spi1_ele1_asyn<5> spi1_n_1930 gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[4] FE_PHN253_SPI_CS spi1_Rx_data_temp<4> spi1_ele1_asyn<4> 
+ FE_PHN263_n_32 spi1_ele1_asyn<4> spi1_n_1930 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[3] FE_PHN253_SPI_CS spi1_Rx_data_temp<3> spi1_ele1_asyn<3> 
+ FE_PHN263_n_32 spi1_ele1_asyn<3> spi1_n_1930 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[2] FE_PHN253_SPI_CS spi1_Rx_data_temp<2> spi1_ele1_asyn<2> 
+ FE_PHN263_n_32 spi1_ele1_asyn<2> spi1_n_1930 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[1] FE_PHN253_SPI_CS spi1_Rx_data_temp<1> spi1_ele1_asyn<1> 
+ FE_PHN263_n_32 spi1_ele1_asyn<1> spi1_n_1930 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_ele1_asyn_reg[0] FE_PHN253_SPI_CS spi1_Rx_data_temp<0> spi1_ele1_asyn<0> 
+ FE_PHN272_FE_OFN33_n_32 spi1_ele1_asyn<0> spi1_n_1930 gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[23] SPI_CS spi1_conf1_asyn<23> spi1_conf1_asyn<23> 
+ FE_PHN431_n_32 spi1_Rx_data_temp<23> spi1_n_1964 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[22] SPI_CS spi1_conf1_asyn<22> spi1_conf1_asyn<22> 
+ FE_PHN431_n_32 spi1_Rx_data_temp<22> spi1_n_1964 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[21] SPI_CS spi1_conf1_asyn<21> spi1_conf1_asyn<21> 
+ FE_PHN431_n_32 spi1_Rx_data_temp<21> spi1_n_1964 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[20] SPI_CS spi1_conf1_asyn<20> spi1_conf1_asyn<20> 
+ FE_PHN431_n_32 spi1_Rx_data_temp<20> spi1_n_1964 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[19] SPI_CS spi1_conf1_asyn<19> spi1_conf1_asyn<19> 
+ FE_PHN431_n_32 spi1_Rx_data_temp<19> spi1_n_1964 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[18] SPI_CS spi1_conf1_asyn<18> spi1_conf1_asyn<18> 
+ FE_PHN431_n_32 spi1_Rx_data_temp<18> spi1_n_1964 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[17] FE_PHN254_SPI_CS spi1_conf1_asyn<17> 
+ spi1_conf1_asyn<17> FE_PHN431_n_32 spi1_Rx_data_temp<17> spi1_n_1964 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[16] FE_PHN254_SPI_CS spi1_conf1_asyn<16> 
+ spi1_conf1_asyn<16> FE_PHN431_n_32 spi1_Rx_data_temp<16> spi1_n_1964 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[15] FE_PHN254_SPI_CS spi1_conf1_asyn<15> 
+ spi1_conf1_asyn<15> FE_PHN431_n_32 spi1_Rx_data_temp<15> spi1_n_1964 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[14] FE_PHN254_SPI_CS spi1_conf1_asyn<14> 
+ spi1_conf1_asyn<14> FE_PHN431_n_32 spi1_Rx_data_temp<14> spi1_n_1964 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[13] FE_PHN254_SPI_CS spi1_conf1_asyn<13> 
+ spi1_conf1_asyn<13> FE_PHN421_n_32 spi1_Rx_data_temp<13> spi1_n_1964 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[12] SPI_CS spi1_conf1_asyn<12> spi1_conf1_asyn<12> 
+ FE_PHN421_n_32 spi1_Rx_data_temp<12> spi1_n_1964 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[11] SPI_CS spi1_conf1_asyn<11> spi1_conf1_asyn<11> 
+ FE_PHN421_n_32 spi1_Rx_data_temp<11> spi1_n_1964 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[10] SPI_CS spi1_conf1_asyn<10> spi1_conf1_asyn<10> 
+ FE_PHN421_n_32 spi1_Rx_data_temp<10> spi1_n_1964 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[9] FE_PHN253_SPI_CS spi1_conf1_asyn<9> spi1_conf1_asyn<9> 
+ FE_OFN443_FE_PHN271_n_32 spi1_Rx_data_temp<9> spi1_n_1964 gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[8] FE_PHN253_SPI_CS spi1_conf1_asyn<8> spi1_conf1_asyn<8> 
+ FE_OFN443_FE_PHN271_n_32 spi1_Rx_data_temp<8> spi1_n_1964 gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[7] FE_PHN253_SPI_CS spi1_conf1_asyn<7> spi1_conf1_asyn<7> 
+ FE_OFN443_FE_PHN271_n_32 spi1_Rx_data_temp<7> spi1_n_1964 gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[6] FE_PHN253_SPI_CS spi1_conf1_asyn<6> spi1_conf1_asyn<6> 
+ FE_OFN443_FE_PHN271_n_32 spi1_Rx_data_temp<6> spi1_n_1964 gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[5] FE_PHN253_SPI_CS spi1_conf1_asyn<5> spi1_conf1_asyn<5> 
+ FE_OFN443_FE_PHN271_n_32 spi1_Rx_data_temp<5> spi1_n_1964 gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[4] FE_PHN253_SPI_CS spi1_conf1_asyn<4> spi1_conf1_asyn<4> 
+ FE_PHN263_n_32 spi1_Rx_data_temp<4> spi1_n_1964 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[3] FE_PHN253_SPI_CS spi1_conf1_asyn<3> spi1_conf1_asyn<3> 
+ FE_PHN263_n_32 spi1_Rx_data_temp<3> spi1_n_1964 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[2] SPI_CS spi1_conf1_asyn<2> spi1_conf1_asyn<2> 
+ FE_PHN421_n_32 spi1_Rx_data_temp<2> spi1_n_1964 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[1] SPI_CS spi1_conf1_asyn<1> spi1_conf1_asyn<1> 
+ FE_PHN263_n_32 spi1_Rx_data_temp<1> spi1_n_1964 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf1_asyn_reg[0] SPI_CS spi1_conf1_asyn<0> spi1_conf1_asyn<0> 
+ FE_PHN421_n_32 spi1_Rx_data_temp<0> spi1_n_1964 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[31] SPI_CS spi1_Rx_data_temp<31> spi1_conf0_asyn<31> 
+ FE_PHN271_n_32 spi1_conf0_asyn<31> spi1_n_2272 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[30] SPI_CS spi1_Rx_data_temp<30> spi1_conf0_asyn<30> 
+ FE_PHN271_n_32 spi1_conf0_asyn<30> spi1_n_2272 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[29] SPI_CS spi1_Rx_data_temp<29> spi1_conf0_asyn<29> 
+ FE_PHN271_n_32 spi1_conf0_asyn<29> spi1_n_2272 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[28] SPI_CS spi1_Rx_data_temp<28> spi1_conf0_asyn<28> 
+ FE_PHN271_n_32 spi1_conf0_asyn<28> spi1_n_2272 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[27] SPI_CS spi1_Rx_data_temp<27> spi1_conf0_asyn<27> 
+ FE_PHN431_n_32 spi1_conf0_asyn<27> spi1_n_2272 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[26] SPI_CS spi1_Rx_data_temp<26> spi1_conf0_asyn<26> 
+ FE_PHN431_n_32 spi1_conf0_asyn<26> spi1_n_2272 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[25] SPI_CS spi1_Rx_data_temp<25> spi1_conf0_asyn<25> 
+ FE_PHN431_n_32 spi1_conf0_asyn<25> spi1_n_2272 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[24] SPI_CS spi1_Rx_data_temp<24> spi1_conf0_asyn<24> 
+ FE_PHN431_n_32 spi1_conf0_asyn<24> spi1_n_2272 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[23] SPI_CS spi1_Rx_data_temp<23> spi1_conf0_asyn<23> 
+ FE_PHN431_n_32 spi1_conf0_asyn<23> spi1_n_2272 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[22] SPI_CS spi1_Rx_data_temp<22> spi1_conf0_asyn<22> 
+ FE_PHN431_n_32 spi1_conf0_asyn<22> spi1_n_2272 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[21] SPI_CS spi1_Rx_data_temp<21> spi1_conf0_asyn<21> 
+ FE_PHN431_n_32 spi1_conf0_asyn<21> spi1_n_2272 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[20] FE_PHN254_SPI_CS spi1_Rx_data_temp<20> 
+ spi1_conf0_asyn<20> FE_PHN421_n_32 spi1_conf0_asyn<20> spi1_n_2272 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[19] SPI_CS spi1_Rx_data_temp<19> spi1_conf0_asyn<19> 
+ FE_OFN33_n_32 spi1_conf0_asyn<19> spi1_n_2272 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[18] SPI_CS spi1_Rx_data_temp<18> spi1_conf0_asyn<18> 
+ FE_PHN421_n_32 spi1_conf0_asyn<18> spi1_n_2272 gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[17] FE_PHN254_SPI_CS spi1_Rx_data_temp<17> 
+ spi1_conf0_asyn<17> FE_PHN421_n_32 spi1_conf0_asyn<17> spi1_n_2272 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[16] FE_PHN254_SPI_CS spi1_Rx_data_temp<16> 
+ spi1_conf0_asyn<16> FE_PHN421_n_32 spi1_conf0_asyn<16> spi1_n_2272 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[15] FE_PHN254_SPI_CS spi1_Rx_data_temp<15> 
+ spi1_conf0_asyn<15> FE_PHN421_n_32 spi1_conf0_asyn<15> spi1_n_2272 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[14] FE_PHN254_SPI_CS spi1_Rx_data_temp<14> 
+ spi1_conf0_asyn<14> FE_PHN421_n_32 spi1_conf0_asyn<14> spi1_n_2272 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[13] FE_PHN254_SPI_CS spi1_Rx_data_temp<13> 
+ spi1_conf0_asyn<13> FE_PHN421_n_32 spi1_conf0_asyn<13> spi1_n_2272 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[12] FE_PHN253_SPI_CS spi1_Rx_data_temp<12> 
+ spi1_conf0_asyn<12> FE_PHN272_FE_OFN33_n_32 spi1_conf0_asyn<12> spi1_n_2272 
+ gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[11] FE_PHN253_SPI_CS spi1_Rx_data_temp<11> 
+ spi1_conf0_asyn<11> FE_OFN443_FE_PHN271_n_32 spi1_conf0_asyn<11> spi1_n_2272 
+ gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[10] FE_PHN253_SPI_CS spi1_Rx_data_temp<10> 
+ spi1_conf0_asyn<10> FE_PHN263_n_32 spi1_conf0_asyn<10> spi1_n_2272 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[9] FE_PHN253_SPI_CS spi1_Rx_data_temp<9> 
+ spi1_conf0_asyn<9> FE_PHN263_n_32 spi1_conf0_asyn<9> spi1_n_2272 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[8] FE_PHN253_SPI_CS spi1_Rx_data_temp<8> 
+ spi1_conf0_asyn<8> FE_PHN263_n_32 spi1_conf0_asyn<8> spi1_n_2272 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[7] FE_PHN253_SPI_CS spi1_Rx_data_temp<7> 
+ spi1_conf0_asyn<7> FE_PHN263_n_32 spi1_conf0_asyn<7> spi1_n_2272 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[6] FE_PHN253_SPI_CS spi1_Rx_data_temp<6> 
+ spi1_conf0_asyn<6> FE_PHN263_n_32 spi1_conf0_asyn<6> spi1_n_2272 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[5] FE_PHN253_SPI_CS spi1_Rx_data_temp<5> 
+ spi1_conf0_asyn<5> FE_PHN263_n_32 spi1_conf0_asyn<5> spi1_n_2272 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[4] FE_PHN253_SPI_CS spi1_Rx_data_temp<4> 
+ spi1_conf0_asyn<4> FE_PHN263_n_32 spi1_conf0_asyn<4> spi1_n_2272 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[3] FE_PHN253_SPI_CS spi1_Rx_data_temp<3> 
+ spi1_conf0_asyn<3> FE_PHN263_n_32 spi1_conf0_asyn<3> spi1_n_2272 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[2] FE_PHN253_SPI_CS spi1_Rx_data_temp<2> 
+ spi1_conf0_asyn<2> FE_PHN263_n_32 spi1_conf0_asyn<2> spi1_n_2272 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[1] FE_PHN253_SPI_CS spi1_Rx_data_temp<1> 
+ spi1_conf0_asyn<1> FE_PHN263_n_32 spi1_conf0_asyn<1> spi1_n_2272 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_conf0_asyn_reg[0] FE_PHN253_SPI_CS spi1_Rx_data_temp<0> 
+ spi1_conf0_asyn<0> FE_PHN263_n_32 spi1_conf0_asyn<0> spi1_n_2272 gnd3i! 
+ vdd3i! / SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[39] CTS_8 spi1_Rx_data_temp<38> spi1_Rx_data_temp<39> 
+ FE_OFN33_n_32 spi1_Rx_data_temp<39> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[38] CTS_8 spi1_Rx_data_temp<37> spi1_Rx_data_temp<38> 
+ FE_OFN33_n_32 spi1_Rx_data_temp<38> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[34] CTS_8 spi1_Rx_data_temp<33> spi1_Rx_data_temp<34> 
+ FE_PHN431_n_32 spi1_Rx_data_temp<34> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[33] CTS_8 spi1_Rx_data_temp<32> spi1_Rx_data_temp<33> 
+ FE_PHN431_n_32 spi1_Rx_data_temp<33> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[32] CTS_8 spi1_Rx_data_temp<31> spi1_Rx_data_temp<32> 
+ FE_PHN431_n_32 spi1_Rx_data_temp<32> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[31] CTS_8 spi1_Rx_data_temp<30> spi1_Rx_data_temp<31> 
+ FE_PHN271_n_32 spi1_Rx_data_temp<31> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[30] CTS_8 spi1_Rx_data_temp<29> spi1_Rx_data_temp<30> 
+ FE_PHN271_n_32 spi1_Rx_data_temp<30> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[29] CTS_8 spi1_Rx_data_temp<28> spi1_Rx_data_temp<29> 
+ FE_PHN271_n_32 spi1_Rx_data_temp<29> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[28] CTS_8 spi1_Rx_data_temp<27> spi1_Rx_data_temp<28> 
+ FE_PHN271_n_32 spi1_Rx_data_temp<28> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[27] CTS_8 spi1_Rx_data_temp<26> spi1_Rx_data_temp<27> 
+ FE_PHN271_n_32 spi1_Rx_data_temp<27> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[26] CTS_8 spi1_Rx_data_temp<25> spi1_Rx_data_temp<26> 
+ FE_PHN271_n_32 spi1_Rx_data_temp<26> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[25] CTS_8 spi1_Rx_data_temp<24> spi1_Rx_data_temp<25> 
+ FE_PHN431_n_32 spi1_Rx_data_temp<25> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[24] CTS_8 spi1_Rx_data_temp<23> spi1_Rx_data_temp<24> 
+ FE_PHN431_n_32 spi1_Rx_data_temp<24> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[23] CTS_8 spi1_Rx_data_temp<22> spi1_Rx_data_temp<23> 
+ FE_OFN35_n_32 spi1_Rx_data_temp<23> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[22] CTS_8 spi1_Rx_data_temp<21> spi1_Rx_data_temp<22> 
+ FE_OFN35_n_32 spi1_Rx_data_temp<22> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[21] CTS_8 spi1_Rx_data_temp<20> spi1_Rx_data_temp<21> 
+ FE_OFN35_n_32 spi1_Rx_data_temp<21> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[20] CTS_8 spi1_Rx_data_temp<19> spi1_Rx_data_temp<20> 
+ FE_OFN35_n_32 spi1_Rx_data_temp<20> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[19] CTS_8 spi1_Rx_data_temp<18> spi1_Rx_data_temp<19> 
+ FE_OFN35_n_32 spi1_Rx_data_temp<19> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[18] CTS_8 spi1_Rx_data_temp<17> spi1_Rx_data_temp<18> 
+ FE_OFN35_n_32 spi1_Rx_data_temp<18> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[17] CTS_8 spi1_Rx_data_temp<16> spi1_Rx_data_temp<17> 
+ FE_PHN431_n_32 spi1_Rx_data_temp<17> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[16] CTS_8 spi1_Rx_data_temp<15> spi1_Rx_data_temp<16> 
+ FE_OFN35_n_32 spi1_Rx_data_temp<16> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[15] CTS_8 spi1_Rx_data_temp<14> spi1_Rx_data_temp<15> 
+ FE_PHN422_n_32 spi1_Rx_data_temp<15> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[14] CTS_8 spi1_Rx_data_temp<13> spi1_Rx_data_temp<14> 
+ FE_PHN422_n_32 spi1_Rx_data_temp<14> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[13] CTS_8 spi1_Rx_data_temp<12> spi1_Rx_data_temp<13> 
+ FE_PHN422_n_32 spi1_Rx_data_temp<13> FE_PHN253_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[12] CTS_8 spi1_Rx_data_temp<11> spi1_Rx_data_temp<12> 
+ FE_PHN422_n_32 spi1_Rx_data_temp<12> FE_PHN253_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[11] CTS_8 spi1_Rx_data_temp<10> spi1_Rx_data_temp<11> 
+ FE_PHN272_FE_OFN33_n_32 spi1_Rx_data_temp<11> FE_PHN253_SPI_CS gnd3i! vdd3i! 
+ / SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[10] CTS_8 spi1_Rx_data_temp<9> spi1_Rx_data_temp<10> 
+ FE_PHN272_FE_OFN33_n_32 spi1_Rx_data_temp<10> FE_PHN253_SPI_CS gnd3i! vdd3i! 
+ / SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[9] CTS_8 spi1_Rx_data_temp<8> spi1_Rx_data_temp<9> 
+ FE_OFN443_FE_PHN271_n_32 spi1_Rx_data_temp<9> FE_PHN253_SPI_CS gnd3i! vdd3i! 
+ / SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[8] CTS_8 spi1_Rx_data_temp<7> spi1_Rx_data_temp<8> 
+ FE_OFN443_FE_PHN271_n_32 spi1_Rx_data_temp<8> FE_PHN253_SPI_CS gnd3i! vdd3i! 
+ / SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[7] CTS_8 spi1_Rx_data_temp<6> spi1_Rx_data_temp<7> 
+ FE_PHN263_n_32 spi1_Rx_data_temp<7> FE_PHN253_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[6] CTS_8 spi1_Rx_data_temp<5> spi1_Rx_data_temp<6> 
+ FE_PHN263_n_32 spi1_Rx_data_temp<6> FE_PHN253_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[5] CTS_8 spi1_Rx_data_temp<4> spi1_Rx_data_temp<5> 
+ FE_PHN263_n_32 spi1_Rx_data_temp<5> FE_PHN253_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[4] CTS_8 spi1_Rx_data_temp<3> spi1_Rx_data_temp<4> 
+ FE_PHN263_n_32 spi1_Rx_data_temp<4> FE_PHN253_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[3] CTS_8 spi1_Rx_data_temp<2> spi1_Rx_data_temp<3> 
+ FE_PHN263_n_32 spi1_Rx_data_temp<3> FE_PHN253_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[2] CTS_8 spi1_Rx_data_temp<1> spi1_Rx_data_temp<2> 
+ FE_PHN263_n_32 spi1_Rx_data_temp<2> FE_PHN253_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[1] CTS_8 spi1_Rx_data_temp<0> spi1_Rx_data_temp<1> 
+ FE_PHN263_n_32 spi1_Rx_data_temp<1> FE_PHN253_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xnpg1_DOWN_count_reg[0] CTS_2 n_356 npg1_DOWN_count<0> FE_PHN422_n_32 n_339 
+ npg1_DOWN_count<0> gnd3i! vdd3i! / SDFRRQJI3VX1
Xnpg1_UP_count_reg[0] CTS_2 n_430 npg1_UP_count<0> FE_PHN422_n_32 n_423 
+ npg1_UP_count<0> gnd3i! vdd3i! / SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[0] CTS_8 FE_PHN274_SPI_MOSI spi1_Rx_data_temp<0> 
+ FE_OFN33_n_32 spi1_Rx_data_temp<0> FE_PHN254_SPI_CS gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[37] CTS_8 spi1_Rx_data_temp<36> spi1_Rx_data_temp<37> 
+ FE_PHN431_n_32 FE_PHN413_spi1_Rx_data_temp_37 FE_PHN254_SPI_CS gnd3i! vdd3i! 
+ / SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[36] CTS_8 spi1_Rx_data_temp<35> spi1_Rx_data_temp<36> 
+ FE_PHN431_n_32 FE_PHN412_spi1_Rx_data_temp_36 FE_PHN254_SPI_CS gnd3i! vdd3i! 
+ / SDFRRQJI3VX1
Xspi1_Rx_data_temp_reg[35] CTS_8 spi1_Rx_data_temp<34> spi1_Rx_data_temp<35> 
+ FE_PHN431_n_32 FE_PHN414_spi1_Rx_data_temp_35 FE_PHN254_SPI_CS gnd3i! vdd3i! 
+ / SDFRRQJI3VX1
Xnpg1_ON_count_reg[0] CTS_2 n_426 npg1_ON_count<0> FE_OFN33_n_32 n_405 
+ npg1_ON_count<0> gnd3i! vdd3i! / SDFRRQJI3VX1
Xnpg1_phase_pause_ready_reg CTS_4 npg1_phase_pause_ready 
+ npg1_phase_pause_ready FE_PHN271_n_32 n_226 n_237 gnd3i! vdd3i! / 
+ SDFRRQJI3VX1
XFE_OFC42_n_510 n_509 FE_OFN40_n_510 gnd3i! vdd3i! / INJI3VX3
Xg9840 npg1_n_374 n_32 gnd3i! vdd3i! / INJI3VX3
XFE_OFC110_enable n_11 enable gnd3i! vdd3i! / INJI3VX3
XFE_OFC121_FE_PHN271_n_32 FE_PHN268_n_32 FE_OFN35_n_32 gnd3i! vdd3i! / INJI3VX3
XFE_OFC123_FE_PHN271_n_32 FE_OFN55_n_32 FE_PHN272_FE_OFN33_n_32 gnd3i! vdd3i! 
+ / INJI3VX3
Xg11813 n_607 up_switches<22> gnd3i! vdd3i! / INJI3VX3
Xg11776 n_612 up_switches<15> gnd3i! vdd3i! / INJI3VX3
Xg11817 n_603 up_switches<14> gnd3i! vdd3i! / INJI3VX3
Xg11742__3680 n_645 n_612 n_603 n_607 n_646 gnd3i! vdd3i! / NA4JI3VX2
Xg11923__5107 npg1_phase_down_state FE_OFN50_npg1_phase_up_state n_510 gnd3i! 
+ vdd3i! / NO2I1JI3VX2
Xg11750__1881 FE_OFN20_up_switches_9 FE_OFN29_up_switches_0 
+ FE_OFN28_up_switches_1 FE_OFN21_up_switches_8 n_638 gnd3i! vdd3i! / OR4JI3VX1
Xg11748__7098 FE_OFN18_up_switches_11 FE_OFN19_up_switches_10 
+ FE_OFN24_up_switches_5 FE_OFN25_up_switches_4 n_640 gnd3i! vdd3i! / OR4JI3VX1
Xg11749__6131 FE_OFN16_up_switches_13 FE_OFN17_up_switches_12 
+ FE_OFN22_up_switches_7 FE_OFN23_up_switches_6 n_639 gnd3i! vdd3i! / OR4JI3VX1
Xg11747__8246 FE_OFN7_up_switches_25 FE_OFN6_up_switches_26 
+ FE_OFN5_up_switches_27 FE_OFN11_up_switches_20 n_641 gnd3i! vdd3i! / 
+ OR4JI3VX1
XFE_OFC94_npg1_phase_up_state FE_OFN50_npg1_phase_up_state 
+ FE_OFN57_npg1_phase_up_state gnd3i! vdd3i! / BUJI3VX2
XFE_OFC44_FE_OFN9_up_switches_23 FE_OFN9_up_switches_23 up_switches<23> gnd3i! 
+ vdd3i! / BUJI3VX2
XFE_OFC41_n_510 n_510 n_509 gnd3i! vdd3i! / BUJI3VX2
XFE_PHC418_SPI_CS FE_PHN415_SPI_CS FE_PHN418_SPI_CS gnd3i! vdd3i! / BUJI3VX2
XFE_OFC153_n_32 FE_PHN422_n_32 FE_PHN263_n_32 gnd3i! vdd3i! / BUJI3VX2
XFE_OFC133_FE_PHN260_n_32 FE_PHN431_n_32 FE_PHN271_n_32 gnd3i! vdd3i! / 
+ BUJI3VX2
XFE_PHC422_n_32 FE_PHN429_n_32 FE_PHN422_n_32 gnd3i! vdd3i! / BUJI3VX2
XFE_OFC45_FE_OFN8_up_switches_24 FE_OFN8_up_switches_24 up_switches<24> gnd3i! 
+ vdd3i! / BUJI3VX2
XFE_OFC43_FE_OFN10_up_switches_21 FE_OFN10_up_switches_21 up_switches<21> 
+ gnd3i! vdd3i! / BUJI3VX2
XFE_PHC413_spi1_Rx_data_temp_37 spi1_Rx_data_temp<37> 
+ FE_PHN413_spi1_Rx_data_temp_37 gnd3i! vdd3i! / BUJI3VX2
XFE_OFC152_n_32 FE_PHN430_n_32 FE_PHN262_n_32 gnd3i! vdd3i! / BUJI3VX2
XCTS_cdb_buf_00030 CTS_6 CTS_3 gnd3i! vdd3i! / BUJI3VX2
XFE_OFC71_FE_OFN14_up_switches_17 FE_OFN14_up_switches_17 up_switches<17> 
+ gnd3i! vdd3i! / BUJI3VX2
XFE_OFC64_FE_OFN15_up_switches_16 FE_OFN15_up_switches_16 up_switches<16> 
+ gnd3i! vdd3i! / BUJI3VX2
XFE_OFC57_FE_OFN1_up_switches_31 FE_OFN1_up_switches_31 up_switches<31> gnd3i! 
+ vdd3i! / BUJI3VX2
XFE_OFC49_FE_OFN2_up_switches_30 FE_OFN2_up_switches_30 up_switches<30> gnd3i! 
+ vdd3i! / BUJI3VX2
XFE_OFC65_FE_OFN4_up_switches_28 FE_OFN4_up_switches_28 up_switches<28> gnd3i! 
+ vdd3i! / BUJI3VX2
XFE_OFC52_FE_OFN3_up_switches_29 FE_OFN3_up_switches_29 up_switches<29> gnd3i! 
+ vdd3i! / BUJI3VX2
XFE_OFC70_FE_OFN12_up_switches_19 FE_OFN12_up_switches_19 up_switches<19> 
+ gnd3i! vdd3i! / BUJI3VX2
XFE_OFC66_FE_OFN13_up_switches_18 FE_OFN13_up_switches_18 up_switches<18> 
+ gnd3i! vdd3i! / BUJI3VX2
XFE_OFC69_FE_OFN6_up_switches_26 FE_OFN6_up_switches_26 up_switches<26> gnd3i! 
+ vdd3i! / BUJI3VX2
XFE_OFC68_FE_OFN7_up_switches_25 FE_OFN7_up_switches_25 up_switches<25> gnd3i! 
+ vdd3i! / BUJI3VX2
XFE_OFC67_FE_OFN5_up_switches_27 FE_OFN5_up_switches_27 up_switches<27> gnd3i! 
+ vdd3i! / BUJI3VX2
XFE_OFC46_FE_OFN11_up_switches_20 FE_OFN11_up_switches_20 up_switches<20> 
+ gnd3i! vdd3i! / BUJI3VX2
XFE_PHC441_n_32 FE_PHN422_n_32 FE_PHN441_n_32 gnd3i! vdd3i! / BUJI3VX3
XFE_PHC433_n_32 FE_PHN422_n_32 FE_PHN433_n_32 gnd3i! vdd3i! / BUJI3VX3
XFE_PHC434_n_32 FE_PHN422_n_32 FE_PHN434_n_32 gnd3i! vdd3i! / BUJI3VX3
XFE_PHC442_n_32 FE_PHN422_n_32 FE_PHN442_n_32 gnd3i! vdd3i! / BUJI3VX3
XFE_PHC436_n_32 FE_PHN422_n_32 FE_PHN436_n_32 gnd3i! vdd3i! / BUJI3VX3
XFE_PHC439_n_32 FE_PHN422_n_32 FE_PHN439_n_32 gnd3i! vdd3i! / BUJI3VX3
XFE_PHC435_n_32 FE_PHN422_n_32 FE_PHN435_n_32 gnd3i! vdd3i! / BUJI3VX3
XFE_PHC430_n_32 FE_PHN421_n_32 FE_PHN430_n_32 gnd3i! vdd3i! / BUJI3VX3
XFE_PHC421_n_32 FE_PHN423_n_32 FE_PHN421_n_32 gnd3i! vdd3i! / BUJI3VX3
XFE_PHC444_n_32 FE_PHN422_n_32 FE_PHN444_n_32 gnd3i! vdd3i! / BUJI3VX3
XFE_PHC443_n_32 FE_PHN422_n_32 FE_PHN443_n_32 gnd3i! vdd3i! / BUJI3VX3
XFE_PHC438_n_32 FE_PHN422_n_32 FE_PHN438_n_32 gnd3i! vdd3i! / BUJI3VX3
XFE_OFC60_FE_OFN28_up_switches_1 FE_OFN28_up_switches_1 up_switches<1> gnd3i! 
+ vdd3i! / BUJI3VX3
XFE_OFC56_FE_OFN20_up_switches_9 FE_OFN20_up_switches_9 up_switches<9> gnd3i! 
+ vdd3i! / BUJI3VX3
XFE_OFC53_FE_OFN21_up_switches_8 FE_OFN21_up_switches_8 up_switches<8> gnd3i! 
+ vdd3i! / BUJI3VX3
XFE_OFC51_FE_OFN29_up_switches_0 FE_OFN29_up_switches_0 up_switches<0> gnd3i! 
+ vdd3i! / BUJI3VX3
XFE_OFC62_FE_OFN27_up_switches_2 FE_OFN27_up_switches_2 up_switches<2> gnd3i! 
+ vdd3i! / BUJI3VX3
XFE_OFC61_FE_OFN26_up_switches_3 FE_OFN26_up_switches_3 up_switches<3> gnd3i! 
+ vdd3i! / BUJI3VX3
XFE_OFC63_FE_OFN25_up_switches_4 FE_OFN25_up_switches_4 up_switches<4> gnd3i! 
+ vdd3i! / BUJI3VX3
XFE_OFC59_FE_OFN24_up_switches_5 FE_OFN24_up_switches_5 up_switches<5> gnd3i! 
+ vdd3i! / BUJI3VX3
XFE_OFC54_FE_OFN19_up_switches_10 FE_OFN19_up_switches_10 up_switches<10> 
+ gnd3i! vdd3i! / BUJI3VX3
XFE_OFC50_FE_OFN18_up_switches_11 FE_OFN18_up_switches_11 up_switches<11> 
+ gnd3i! vdd3i! / BUJI3VX3
XFE_OFC58_FE_OFN23_up_switches_6 FE_OFN23_up_switches_6 up_switches<6> gnd3i! 
+ vdd3i! / BUJI3VX3
XFE_OFC55_FE_OFN22_up_switches_7 FE_OFN22_up_switches_7 up_switches<7> gnd3i! 
+ vdd3i! / BUJI3VX3
XFE_OFC48_FE_OFN17_up_switches_12 FE_OFN17_up_switches_12 up_switches<12> 
+ gnd3i! vdd3i! / BUJI3VX3
XFE_OFC47_FE_OFN16_up_switches_13 FE_OFN16_up_switches_13 up_switches<13> 
+ gnd3i! vdd3i! / BUJI3VX3
Xg11780__2883 FE_OFN40_n_510 n_514 n_600 down_switches<2> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11832__2802 FE_OFN40_n_510 n_536 n_599 down_switches<8> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11825__6260 FE_OFN40_n_510 n_522 n_597 down_switches<6> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11779__9945 FE_OFN40_n_510 n_520 n_596 down_switches<3> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11833__1705 FE_OFN40_n_510 n_540 n_594 down_switches<17> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11781__2346 FE_OFN40_n_510 n_535 n_593 down_switches<1> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11836__7098 FE_OFN40_n_510 n_526 n_592 down_switches<9> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11782__1666 FE_OFN40_n_510 n_530 n_591 down_switches<0> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11830__3680 FE_OFN40_n_510 n_543 n_588 down_switches<19> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11783__7410 FE_OFN40_n_510 n_534 n_582 down_switches<31> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11827__8428 FE_OFN40_n_510 n_532 n_579 down_switches<21> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11826__4319 FE_OFN40_n_510 n_529 n_574 down_switches<22> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11828__5526 FE_OFN40_n_510 n_518 n_572 down_switches<7> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11778__9315 FE_OFN40_n_510 n_517 n_569 down_switches<28> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11824__5107 FE_OFN40_n_510 n_515 n_567 down_switches<23> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11837__6131 FE_OFN40_n_510 n_516 n_566 down_switches<10> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11831__1617 FE_OFN40_n_510 n_523 n_565 down_switches<18> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11821__6417 FE_OFN40_n_510 n_521 n_564 down_switches<5> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11841__4733 FE_OFN40_n_510 n_525 n_563 down_switches<11> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11822__5477 FE_OFN40_n_510 n_539 n_562 down_switches<25> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11823__2398 FE_OFN40_n_510 n_528 n_560 down_switches<24> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11820__7410 FE_OFN40_n_510 n_541 n_559 down_switches<26> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11784__6417 FE_OFN40_n_510 n_519 n_558 down_switches<30> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11829__6783 FE_OFN40_n_510 n_538 n_556 down_switches<20> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11835__8246 FE_OFN40_n_510 n_524 n_555 down_switches<27> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11785__5477 FE_OFN40_n_510 n_533 n_554 down_switches<29> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11786__2398 FE_OFN40_n_510 n_542 n_553 down_switches<4> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11834__5122 FE_OFN40_n_510 n_513 n_552 down_switches<16> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11840__7482 FE_OFN40_n_510 n_531 n_549 down_switches<12> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11839__5115 FE_OFN40_n_510 n_544 n_548 down_switches<13> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11838__1881 FE_OFN40_n_510 n_537 n_547 down_switches<14> gnd3i! vdd3i! / 
+ ON21JI3VX4
Xg11819__1666 FE_OFN40_n_510 n_527 n_545 down_switches<15> gnd3i! vdd3i! / 
+ ON21JI3VX4
XFE_PHC254_SPI_CS FE_PHN418_SPI_CS FE_PHN254_SPI_CS gnd3i! vdd3i! / BUJI3VX1
XFE_OFC157_FE_PHN254_SPI_CS FE_PHN254_SPI_CS FE_PHN253_SPI_CS gnd3i! vdd3i! / 
+ BUJI3VX1
XCTS_cdb_buf_00028 CTS_10 CTS_9 gnd3i! vdd3i! / BUJI3VX1
XCTS_cdb_buf_00027 CTS_11 CTS_10 gnd3i! vdd3i! / BUJI3VX1
XCTS_cdb_buf_00026 SPI_Clk CTS_11 gnd3i! vdd3i! / BUJI3VX1
XFE_PHC428_n_32 FE_PHN430_n_32 FE_PHN428_n_32 gnd3i! vdd3i! / BUJI3VX1
XFE_PHC427_n_32 FE_PHN448_n_32 FE_PHN427_n_32 gnd3i! vdd3i! / BUJI3VX1
XCTS_cdb_buf_00032 CTS_7 CTS_6 gnd3i! vdd3i! / BUJI3VX1
XCTS_cdb_buf_00031 clk CTS_7 gnd3i! vdd3i! / BUJI3VX1
XFE_OFC108_npg1_phase_down_state npg1_phase_down_state 
+ FE_OFN58_npg1_phase_down_state gnd3i! vdd3i! / BUJI3VX1
XFE_OFC156_FE_PHN254_SPI_CS FE_PHN254_SPI_CS FE_OFN30_SPI_CS gnd3i! vdd3i! / 
+ INJI3VX1
XFE_OFC122_FE_PHN271_n_32 FE_PHN268_n_32 FE_OFN33_n_32 gnd3i! vdd3i! / INJI3VX1
XFE_OFC150_n_32 FE_PHN422_n_32 FE_PHN268_n_32 gnd3i! vdd3i! / INJI3VX1
XFE_OFC151_n_32 FE_PHN422_n_32 FE_OFN55_n_32 gnd3i! vdd3i! / INJI3VX1
XFE_OFC160_npg1_OFF_count_3 npg1_OFF_count<3> FE_PHN233_npg1_OFF_count_3 
+ gnd3i! vdd3i! / INJI3VX1
XFE_OFC159_npg1_OFF_count_0 npg1_OFF_count<0> n_44 gnd3i! vdd3i! / INJI3VX1
XFE_OFC109_enable FE_OFN52_enable n_11 gnd3i! vdd3i! / INJI3VX1
XFE_OFC164_npg1_phase_down_count_1 npg1_phase_down_count<1> n_22 gnd3i! vdd3i! 
+ / INJI3VX1
XFE_OFC163_npg1_freq_count_6 npg1_freq_count<6> n_43 gnd3i! vdd3i! / INJI3VX1
XFE_OFC162_npg1_freq_count_5 npg1_freq_count<5> n_52 gnd3i! vdd3i! / INJI3VX1
XFE_OFC161_npg1_freq_count_3 npg1_freq_count<3> n_42 gnd3i! vdd3i! / INJI3VX1
XFE_OFC158_npg1_freq_count_10 npg1_freq_count<10> n_54 gnd3i! vdd3i! / INJI3VX1
XFE_OFC124_FE_PHN271_n_32 FE_OFN55_n_32 FE_OFN443_FE_PHN271_n_32 gnd3i! vdd3i! 
+ / INJI3VX2
Xg17164 n_736 ele1<16> FE_OFN15_up_switches_16 FE_OFN50_npg1_phase_up_state 
+ gnd3i! vdd3i! / MU2JI3VX0
Xg17162 n_734 ele1<31> FE_OFN1_up_switches_31 FE_OFN50_npg1_phase_up_state 
+ gnd3i! vdd3i! / MU2JI3VX0
Xg17160 n_732 ele1<30> FE_OFN2_up_switches_30 FE_OFN50_npg1_phase_up_state 
+ gnd3i! vdd3i! / MU2JI3VX0
Xg2 n_730 ele1<29> FE_OFN3_up_switches_29 FE_OFN50_npg1_phase_up_state gnd3i! 
+ vdd3i! / MU2JI3VX0
XCTS_cdb_buf_00025 CTS_9 CTS_8 gnd3i! vdd3i! / BUJI3VX6
XFE_PHC431_n_32 FE_PHN262_n_32 FE_PHN431_n_32 gnd3i! vdd3i! / BUJI3VX6
XFE_OFC99_pulse_active FE_OFN39_pulse_active pulse_active gnd3i! vdd3i! / 
+ BUJI3VX6
XFE_OFC93_npg1_phase_up_state npg1_phase_up_state FE_OFN50_npg1_phase_up_state 
+ gnd3i! vdd3i! / BUJI3VX6
Xg11743__1617 n_644 n_641 n_642 n_645 gnd3i! vdd3i! / NO3JI3VX1
Xg11741__6783 n_646 n_639 n_643 n_640 FE_OFN39_pulse_active gnd3i! vdd3i! / 
+ OR4JI3VX2
Xg16582__3680 n_497 npg1_UP_accumulator<9> conf1<9> n_501 gnd3i! vdd3i! / 
+ EO3JI3VX1
Xg16581__6783 n_499 npg1_DOWN_accumulator<9> conf1<9> n_502 gnd3i! vdd3i! / 
+ EO3JI3VX1
XFE_PHC415_SPI_CS FE_PHN275_SPI_CS FE_PHN415_SPI_CS gnd3i! vdd3i! / BUJI3VX16
XFE_PHC447_n_32 FE_PHN422_n_32 FE_PHN447_n_32 gnd3i! vdd3i! / BUJI3VX16
XFE_PHC446_n_32 FE_PHN422_n_32 FE_PHN446_n_32 gnd3i! vdd3i! / BUJI3VX16
XFE_PHC445_n_32 FE_PHN422_n_32 FE_PHN445_n_32 gnd3i! vdd3i! / BUJI3VX16
XFE_PHC274_SPI_MOSI FE_PHN416_SPI_MOSI FE_PHN274_SPI_MOSI gnd3i! vdd3i! / 
+ DLY4JI3VX1
Xspi1_Rx_count_reg[2] CTS_8 spi1_n_1999 spi1_Rx_count<2> FE_OFN30_SPI_CS 
+ gnd3i! vdd3i! / DFRRQJI3VX2
XFE_PHC440_n_32 FE_PHN422_n_32 FE_PHN440_n_32 gnd3i! vdd3i! / DLY2JI3VX1
Xspi1_g2__6417 spi1_n_1994 spi1_Rx_data_temp<33> spi1_n_2271 gnd3i! vdd3i! / 
+ NA2I1JI3VX2
Xspi1_g996__5477 spi1_Rx_data_temp<33> spi1_n_1995 spi1_n_2272 gnd3i! vdd3i! / 
+ NA2I1JI3VX2
Xspi1_g934__7098 spi1_n_1995 spi1_Rx_data_temp<33> spi1_n_1930 gnd3i! vdd3i! / 
+ NA2JI3VX2
Xspi1_g936__6131 spi1_n_1994 spi1_Rx_data_temp<33> spi1_n_1964 gnd3i! vdd3i! / 
+ NO2JI3VX2
XFILLCAP_T_1_6 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_7 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_12 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_19 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_22 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_24 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_26 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_38 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_39 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_40 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_44 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_45 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_51 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_59 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_63 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_64 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_72 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_73 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_75 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_80 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_87 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_96 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_103 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_104 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_105 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_107 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_108 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_111 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_118 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_120 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_121 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_123 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_125 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_132 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_133 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_134 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_136 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_137 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_140 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_141 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_150 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_158 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_159 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_160 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_164 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_165 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_185 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_194 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_197 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_199 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_212 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_219 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_226 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_229 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_231 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_233 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_254 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_260 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_265 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_272 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_276 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_280 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_283 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_306 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_311 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_314 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_319 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_344 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_347 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_355 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_363 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_364 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_366 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_373 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_378 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_379 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_387 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_389 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_390 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_400 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_403 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_405 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_409 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_414 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_415 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_420 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_421 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_440 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_444 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_445 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_450 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_452 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_453 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_462 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_467 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_468 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_469 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_471 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_474 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_475 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_484 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_493 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_498 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_501 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_502 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_507 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_511 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_514 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_521 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_523 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_528 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_530 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_532 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_534 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_537 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_552 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_553 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_555 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_560 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_563 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_569 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_576 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_584 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_597 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_608 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_609 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_632 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_638 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_648 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_657 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_667 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_690 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_705 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_707 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_710 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_711 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_719 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_727 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_730 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_741 gnd3i! vdd3i! / DECAP5JI3V
XFILLCAP_T_1_3 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_4 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_5 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_8 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_11 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_15 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_16 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_17 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_18 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_20 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_21 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_23 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_28 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_29 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_30 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_33 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_34 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_35 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_36 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_37 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_42 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_43 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_47 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_48 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_49 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_50 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_53 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_54 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_55 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_56 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_57 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_58 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_60 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_61 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_67 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_68 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_70 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_71 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_74 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_78 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_82 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_83 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_85 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_86 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_88 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_89 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_91 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_92 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_94 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_98 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_99 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_101 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_102 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_109 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_113 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_114 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_116 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_117 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_119 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_124 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_126 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_128 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_129 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_135 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_138 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_139 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_144 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_145 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_149 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_151 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_152 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_153 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_154 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_155 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_156 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_157 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_161 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_162 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_167 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_168 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_170 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_171 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_172 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_174 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_175 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_176 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_177 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_178 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_179 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_180 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_181 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_182 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_183 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_187 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_188 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_193 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_195 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_201 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_202 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_206 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_207 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_208 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_210 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_211 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_214 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_215 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_216 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_217 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_218 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_222 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_223 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_224 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_225 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_228 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_235 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_236 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_237 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_239 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_241 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_242 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_245 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_247 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_248 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_249 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_250 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_253 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_259 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_262 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_263 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_264 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_267 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_268 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_269 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_270 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_271 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_278 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_279 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_281 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_282 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_285 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_286 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_287 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_288 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_289 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_290 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_292 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_293 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_295 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_296 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_298 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_299 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_300 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_301 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_305 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_308 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_309 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_310 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_313 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_315 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_316 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_317 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_318 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_321 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_325 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_327 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_328 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_329 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_330 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_331 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_333 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_334 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_335 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_337 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_338 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_339 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_340 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_343 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_345 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_348 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_351 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_352 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_356 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_357 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_358 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_359 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_361 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_362 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_368 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_375 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_376 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_377 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_380 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_381 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_382 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_383 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_384 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_385 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_386 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_394 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_395 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_397 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_398 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_399 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_402 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_408 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_417 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_418 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_419 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_423 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_424 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_425 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_426 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_428 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_429 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_434 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_435 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_437 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_438 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_439 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_442 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_443 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_448 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_449 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_455 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_456 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_458 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_459 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_460 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_461 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_464 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_465 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_466 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_470 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_477 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_478 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_479 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_482 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_483 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_485 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_491 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_492 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_496 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_497 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_503 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_504 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_505 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_513 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_518 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_520 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_526 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_533 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_539 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_540 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_542 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_545 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_546 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_547 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_548 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_549 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_551 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_554 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_556 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_559 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_561 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_564 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_565 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_566 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_567 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_568 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_570 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_574 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_575 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_578 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_579 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_582 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_583 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_585 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_586 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_587 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_591 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_592 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_593 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_595 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_598 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_600 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_601 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_606 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_610 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_611 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_618 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_620 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_621 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_622 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_623 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_624 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_625 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_634 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_636 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_639 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_640 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_645 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_646 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_647 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_651 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_652 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_653 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_654 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_655 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_663 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_664 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_669 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_670 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_671 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_672 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_673 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_674 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_681 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_684 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_685 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_686 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_687 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_688 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_689 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_701 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_702 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_703 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_704 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_708 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_718 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_723 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_724 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_725 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_726 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_728 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_729 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_737 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_738 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_739 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_740 gnd3i! vdd3i! / DECAP7JI3V
XFILLCAP_T_1_2 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_10 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_25 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_46 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_52 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_62 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_65 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_90 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_93 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_97 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_106 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_110 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_112 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_127 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_131 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_142 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_148 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_173 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_190 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_191 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_192 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_196 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_198 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_204 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_205 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_209 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_213 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_220 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_221 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_230 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_232 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_234 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_240 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_261 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_297 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_302 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_307 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_312 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_320 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_323 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_324 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_332 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_336 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_349 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_350 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_354 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_388 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_391 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_404 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_407 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_411 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_416 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_422 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_431 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_441 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_447 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_463 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_473 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_488 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_489 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_495 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_506 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_510 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_517 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_519 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_525 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_529 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_541 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_550 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_605 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_607 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_612 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_614 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_626 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_635 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_637 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_644 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_658 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_680 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_683 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_691 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_700 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_706 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_709 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_717 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_731 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_736 gnd3i! vdd3i! / DECAP15JI3V
XFILLCAP_T_1_1 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_9 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_13 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_27 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_31 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_32 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_69 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_81 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_84 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_100 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_115 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_130 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_146 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_147 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_166 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_169 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_186 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_189 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_200 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_203 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_227 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_243 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_251 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_252 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_255 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_257 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_266 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_273 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_274 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_275 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_277 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_294 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_303 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_322 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_341 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_342 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_346 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_353 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_360 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_365 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_370 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_374 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_392 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_396 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_406 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_410 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_412 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_413 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_430 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_451 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_454 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_472 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_476 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_486 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_487 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_494 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_499 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_508 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_509 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_515 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_516 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_524 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_535 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_536 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_543 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_557 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_558 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_572 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_588 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_589 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_590 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_602 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_603 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_604 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_615 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_616 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_617 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_628 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_629 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_630 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_631 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_641 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_642 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_643 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_649 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_656 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_659 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_660 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_661 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_662 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_665 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_666 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_675 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_676 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_677 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_678 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_679 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_682 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_692 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_693 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_694 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_695 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_696 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_697 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_698 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_699 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_712 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_713 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_714 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_715 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_716 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_720 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_721 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_722 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_732 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_733 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_734 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_735 gnd3i! vdd3i! / DECAP25JI3V
XFILLCAP_T_1_14 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_41 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_66 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_76 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_77 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_79 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_95 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_122 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_143 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_163 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_184 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_238 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_244 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_246 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_256 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_258 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_284 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_291 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_304 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_326 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_367 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_369 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_371 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_372 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_393 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_401 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_427 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_432 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_433 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_436 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_446 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_457 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_480 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_481 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_490 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_500 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_512 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_522 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_527 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_531 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_538 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_544 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_562 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_571 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_573 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_577 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_580 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_581 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_594 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_596 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_599 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_613 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_619 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_627 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_633 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_650 gnd3i! vdd3i! / DECAP10JI3V
XFILLCAP_T_1_668 gnd3i! vdd3i! / DECAP10JI3V
.ENDS

