* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : aska_dig_lvs                                 *
* Netlisted  : Mon Sep  9 14:36:59 2024                     *
* PVS Version: 23.10-p043 Mon Oct 2 18:09:08 PDT 2023      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(ne3i) nemi ndiff(D) p1trm(G) ndiff(S) pwitrm(B)
*.DEVTMPLT 1 MP(pe3i) pemi pdiff(D) p1trm(G) pdiff(S) dnwtrm(B)
*.DEVTMPLT 2 D(p_ddnwmv) p_ddnwmv bulk(POS) dnwtrm(NEG)
*.DEVTMPLT 3 D(p_dipdnwmv) p_dipwmv pwitrm(POS) dnwtrm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: EN2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt EN2JI3VX0 vdd3i! gnd3i! A B Q
*.DEVICECLIMB
** N=10 EP=5 FDC=10
M0 8 A 9 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=620 $Y=980 $dt=0
M1 gnd3i! B 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=1220 $Y=980 $dt=0
M2 7 A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=1.134e-13 PD=9.6e-07 PS=9.6e-07 $X=2110 $Y=980 $dt=0
M3 gnd3i! B 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.698e-13 AS=1.134e-13 PD=3.22e-06 PS=9.6e-07 $X=3000 $Y=980 $dt=0
M4 Q 9 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=2.058e-13 PD=1.8e-06 PS=1.82e-06 $X=4440 $Y=1020 $dt=0
M5 9 A vdd3i! vdd3i! pe3i L=3e-07 W=9e-07 AD=3.195e-13 AS=8.517e-13 PD=1.61e-06 PS=4.61e-06 $X=685 $Y=2410 $dt=1
M6 vdd3i! B 9 vdd3i! pe3i L=3e-07 W=9e-07 AD=4.30855e-13 AS=3.195e-13 PD=1.83273e-06 PS=1.61e-06 $X=1695 $Y=2410 $dt=1
M7 10 A vdd3i! vdd3i! pe3i L=3e-07 W=1.3e-06 AD=1.95e-13 AS=6.22345e-13 PD=1.6e-06 PS=2.64727e-06 $X=2825 $Y=2520 $dt=1
M8 Q B 10 vdd3i! pe3i L=3e-07 W=1.3e-06 AD=6.21324e-13 AS=1.95e-13 PD=2.52941e-06 PS=1.6e-06 $X=3425 $Y=2520 $dt=1
M9 vdd3i! 9 Q vdd3i! pe3i L=3e-07 W=9.1e-07 AD=8.0675e-13 AS=4.34926e-13 PD=4.39e-06 PS=1.77059e-06 $X=4575 $Y=2520 $dt=1
.ends EN2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO3JI3VX1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO3JI3VX1 vdd3i! gnd3i! C Q B A
*.DEVICECLIMB
** N=9 EP=6 FDC=6
M0 Q C gnd3i! gnd3i! ne3i L=3.4986e-07 W=8.92071e-07 AD=2.37813e-13 AS=4.30337e-13 PD=1.42707e-06 PS=2.76707e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! B Q gnd3i! ne3i L=3.4986e-07 W=8.92071e-07 AD=2.40287e-13 AS=2.37813e-13 PD=1.44207e-06 PS=1.42707e-06 $X=1500 $Y=660 $dt=0
M2 Q A gnd3i! gnd3i! ne3i L=3.4986e-07 W=8.92071e-07 AD=4.29162e-13 AS=2.40287e-13 PD=2.74707e-06 PS=1.44207e-06 $X=2390 $Y=660 $dt=0
M3 9 C vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=1.3994e-12 PD=1.72e-06 PS=5.15e-06 $X=955 $Y=2410 $dt=1
M4 8 B 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=2.1855e-13 PD=1.72e-06 PS=1.72e-06 $X=1565 $Y=2410 $dt=1
M5 Q A 8 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=2.1855e-13 PD=3.78e-06 PS=1.72e-06 $X=2175 $Y=2410 $dt=1
.ends NO3JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA2JI3VX2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA2JI3VX2 vdd3i! gnd3i! B Q A
*.DEVICECLIMB
** N=8 EP=5 FDC=8
M0 8 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=7.09e-13 PD=1.14e-06 PS=3.68e-06 $X=740 $Y=660 $dt=0
M1 Q A 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=1.1125e-13 PD=1.43e-06 PS=1.14e-06 $X=1340 $Y=660 $dt=0
M2 7 A Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=2.403e-13 PD=1.14e-06 PS=1.43e-06 $X=2230 $Y=660 $dt=0
M3 gnd3i! B 7 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=7.09e-13 AS=1.1125e-13 PD=3.68e-06 PS=1.14e-06 $X=2830 $Y=660 $dt=0
M4 Q B vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.7e-13 AS=8.172e-13 PD=1.54e-06 PS=4.22e-06 $X=540 $Y=2410 $dt=1
M5 vdd3i! A Q vdd3i! pe3i L=3e-07 W=1e-06 AD=8.172e-13 AS=2.7e-13 PD=4.22e-06 PS=1.54e-06 $X=1380 $Y=2410 $dt=1
M6 Q A vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.7e-13 AS=8.172e-13 PD=1.54e-06 PS=4.22e-06 $X=2240 $Y=2410 $dt=1
M7 vdd3i! B Q vdd3i! pe3i L=3e-07 W=1e-06 AD=8.172e-13 AS=2.7e-13 PD=4.22e-06 PS=1.54e-06 $X=3080 $Y=2410 $dt=1
.ends NA2JI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO22JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO22JI3VX1 vdd3i! gnd3i! B A Q C
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 8 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=4.87734e-13 PD=9.6e-07 PS=2.24324e-06 $X=720 $Y=1130 $dt=0
M1 gnd3i! A 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=4.87734e-13 AS=1.134e-13 PD=2.24324e-06 PS=9.6e-07 $X=1610 $Y=1130 $dt=0
M2 Q 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=1.03353e-12 PD=1.43e-06 PS=4.75353e-06 $X=2580 $Y=660 $dt=0
M3 gnd3i! C Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=6.098e-13 AS=2.403e-13 PD=3.52e-06 PS=1.43e-06 $X=3470 $Y=660 $dt=0
M4 10 B vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=1.0178e-12 PD=1.1e-06 PS=4.78e-06 $X=770 $Y=2410 $dt=1
M5 8 A 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.505e-13 AS=1.0625e-13 PD=2.76e-06 PS=1.1e-06 $X=1320 $Y=2410 $dt=1
M6 9 8 Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=6.768e-13 PD=1.66e-06 PS=3.78e-06 $X=2920 $Y=2410 $dt=1
M7 vdd3i! C 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=9.682e-13 AS=1.7625e-13 PD=4.66e-06 PS=1.66e-06 $X=3470 $Y=2410 $dt=1
.ends NO22JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DFRRQJI3VX2                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DFRRQJI3VX2 vdd3i! gnd3i! RN D C Q
*.DEVICECLIMB
** N=23 EP=6 FDC=32
M0 gnd3i! 17 19 gnd3i! ne3i L=3.5e-07 W=6.6e-07 AD=1.94849e-13 AS=3.168e-13 PD=1.21781e-06 PS=2.28e-06 $X=620 $Y=660 $dt=0
M1 10 RN gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.28952e-13 AS=2.62751e-13 PD=2.36956e-06 PS=1.64219e-06 $X=1510 $Y=660 $dt=0
M2 18 19 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.55236e-13 PD=6.7e-07 PS=1.11822e-06 $X=2340 $Y=1390 $dt=0
M3 17 9 18 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=2940 $Y=1390 $dt=0
M4 16 15 17 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=3830 $Y=1390 $dt=0
M5 10 D 16 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.835e-13 AS=5.25e-14 PD=2.19e-06 PS=6.7e-07 $X=4430 $Y=1390 $dt=0
M6 gnd3i! C 15 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.659e-13 AS=2.016e-13 PD=1.21e-06 PS=1.8e-06 $X=6060 $Y=1390 $dt=0
M7 9 15 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.95e-13 AS=1.659e-13 PD=2.23e-06 PS=1.21e-06 $X=7045 $Y=1390 $dt=0
M8 14 19 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=8695 $Y=1020 $dt=0
M9 13 9 14 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=9295 $Y=1020 $dt=0
M10 12 15 13 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=10185 $Y=1020 $dt=0
M11 8 11 12 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.55817e-13 AS=5.25e-14 PD=9.68244e-07 PS=6.7e-07 $X=10785 $Y=1020 $dt=0
M12 gnd3i! RN 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=5.94987e-13 AS=3.30183e-13 PD=3.35209e-06 PS=2.05176e-06 $X=11755 $Y=660 $dt=0
M13 11 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=6.6e-07 AD=3.168e-13 AS=4.41226e-13 PD=2.28e-06 PS=2.48582e-06 $X=12750 $Y=890 $dt=0
M14 Q 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=5.94987e-13 PD=1.43e-06 PS=3.35209e-06 $X=14380 $Y=660 $dt=0
M15 gnd3i! 13 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=2.403e-13 PD=2.74e-06 PS=1.43e-06 $X=15270 $Y=660 $dt=0
M16 vdd3i! 17 19 vdd3i! pe3i L=3e-07 W=1e-06 AD=2.97674e-13 AS=4.8e-13 PD=1.7907e-06 PS=2.96e-06 $X=620 $Y=2670 $dt=1
M17 17 RN vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.136e-13 AS=2.14326e-13 PD=2.4e-06 PS=1.2893e-06 $X=1460 $Y=2670 $dt=1
M18 23 19 vdd3i! vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=5.1875e-13 PD=6.7e-07 PS=2.99e-06 $X=3080 $Y=3400 $dt=1
M19 17 15 23 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=1.21617e-13 AS=5.25e-14 PD=9.13043e-07 PS=6.7e-07 $X=3630 $Y=3400 $dt=1
M20 22 9 17 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=1.2e-13 AS=2.77983e-13 PD=1.21e-06 PS=2.08696e-06 $X=4470 $Y=2860 $dt=1
M21 vdd3i! D 22 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=5.00229e-13 AS=1.2e-13 PD=2.34286e-06 PS=1.21e-06 $X=5020 $Y=2860 $dt=1
M22 15 C vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=4.56625e-13 AS=3.75171e-13 PD=2.86e-06 PS=1.75714e-06 $X=6060 $Y=2860 $dt=1
M23 vdd3i! 15 9 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.92547e-13 AS=3.528e-13 PD=1.8586e-06 PS=2.42e-06 $X=7720 $Y=2670 $dt=1
M24 21 19 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=1.25e-13 AS=5.45203e-13 PD=1.25e-06 PS=2.5814e-06 $X=8740 $Y=2820 $dt=1
M25 13 15 21 vdd3i! pe3i L=3e-07 W=1e-06 AD=2.96338e-13 AS=1.25e-13 PD=2.19718e-06 PS=1.25e-06 $X=9290 $Y=2820 $dt=1
M26 20 9 13 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=1.24462e-13 PD=6.7e-07 PS=9.22817e-07 $X=10150 $Y=3235 $dt=1
M27 vdd3i! 11 20 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=3.93439e-13 AS=5.25e-14 PD=1.64096e-06 PS=6.7e-07 $X=10700 $Y=3235 $dt=1
M28 vdd3i! RN 13 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=6.74468e-13 AS=2.976e-13 PD=2.81307e-06 PS=2.4e-06 $X=11900 $Y=2410 $dt=1
M29 11 13 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=4.8e-13 AS=9.36761e-13 PD=2.96e-06 PS=3.90704e-06 $X=12740 $Y=2410 $dt=1
M30 Q 13 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=1.32083e-12 PD=1.95e-06 PS=5.50893e-06 $X=14440 $Y=2410 $dt=1
M31 vdd3i! 13 Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=8.802e-13 AS=3.807e-13 PD=4.56e-06 PS=1.95e-06 $X=15280 $Y=2410 $dt=1
.ends DFRRQJI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX8                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX8 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=19
M0 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=6.098e-13 PD=1.43e-06 PS=3.52e-06 $X=660 $Y=660 $dt=0
M1 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.804e-13 AS=2.403e-13 PD=1.91e-06 PS=1.43e-06 $X=1550 $Y=660 $dt=0
M2 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.804e-13 PD=1.43e-06 PS=1.91e-06 $X=2570 $Y=660 $dt=0
M3 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=3460 $Y=660 $dt=0
M4 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=4430 $Y=660 $dt=0
M5 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=5320 $Y=660 $dt=0
M6 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=6290 $Y=660 $dt=0
M7 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=8.702e-13 AS=2.403e-13 PD=3.94e-06 PS=1.43e-06 $X=7180 $Y=660 $dt=0
M8 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=5.51013e-13 PD=1.86506e-06 PS=3.69506e-06 $X=620 $Y=2410 $dt=1
M9 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.61963e-13 AS=2.83187e-13 PD=1.87506e-06 PS=1.86506e-06 $X=1170 $Y=2410 $dt=1
M10 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.61963e-13 PD=1.86506e-06 PS=1.87506e-06 $X=2020 $Y=2410 $dt=1
M11 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.61963e-13 AS=2.83187e-13 PD=1.87506e-06 PS=1.86506e-06 $X=2570 $Y=2410 $dt=1
M12 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.61963e-13 PD=1.86506e-06 PS=1.87506e-06 $X=3420 $Y=2410 $dt=1
M13 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.61963e-13 AS=2.83187e-13 PD=1.87506e-06 PS=1.86506e-06 $X=3970 $Y=2410 $dt=1
M14 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.61963e-13 PD=1.86506e-06 PS=1.87506e-06 $X=4820 $Y=2410 $dt=1
M15 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.61963e-13 AS=2.83187e-13 PD=1.87506e-06 PS=1.86506e-06 $X=5370 $Y=2410 $dt=1
M16 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.61963e-13 PD=1.86506e-06 PS=1.87506e-06 $X=6220 $Y=2410 $dt=1
M17 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.61963e-13 AS=2.83187e-13 PD=1.87506e-06 PS=1.86506e-06 $X=6770 $Y=2410 $dt=1
M18 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=5.79287e-13 AS=2.61963e-13 PD=3.69506e-06 PS=1.87506e-06 $X=7620 $Y=2410 $dt=1
.ends BUJI3VX8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DFRRQJI3VX4                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DFRRQJI3VX4 vdd3i! gnd3i! RN D C Q
*.DEVICECLIMB
** N=23 EP=6 FDC=36
M0 gnd3i! 17 19 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=4.272e-13 PD=1.43e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 10 RN gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.28952e-13 AS=2.403e-13 PD=2.36956e-06 PS=1.43e-06 $X=1510 $Y=660 $dt=0
M2 18 19 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.55236e-13 PD=6.7e-07 PS=1.11822e-06 $X=2340 $Y=1390 $dt=0
M3 17 9 18 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=2940 $Y=1390 $dt=0
M4 16 15 17 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=3830 $Y=1390 $dt=0
M5 10 D 16 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.835e-13 AS=5.25e-14 PD=2.19e-06 PS=6.7e-07 $X=4430 $Y=1390 $dt=0
M6 gnd3i! C 15 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.659e-13 AS=2.016e-13 PD=1.21e-06 PS=1.8e-06 $X=6060 $Y=1390 $dt=0
M7 9 15 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.95e-13 AS=1.659e-13 PD=2.23e-06 PS=1.21e-06 $X=7045 $Y=1390 $dt=0
M8 14 19 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=8695 $Y=1020 $dt=0
M9 13 9 14 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=9295 $Y=1020 $dt=0
M10 12 15 13 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=10185 $Y=1020 $dt=0
M11 8 11 12 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.55817e-13 AS=5.25e-14 PD=9.68244e-07 PS=6.7e-07 $X=10785 $Y=1020 $dt=0
M12 gnd3i! RN 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.60325e-13 AS=3.30183e-13 PD=1.475e-06 PS=2.05176e-06 $X=11755 $Y=660 $dt=0
M13 11 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=2.60325e-13 PD=2.74e-06 PS=1.475e-06 $X=12690 $Y=660 $dt=0
M14 Q 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=4.272e-13 PD=1.43e-06 PS=2.74e-06 $X=14280 $Y=660 $dt=0
M15 gnd3i! 13 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=15170 $Y=660 $dt=0
M16 Q 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=16060 $Y=660 $dt=0
M17 gnd3i! 13 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=2.403e-13 PD=2.74e-06 PS=1.43e-06 $X=16950 $Y=660 $dt=0
M18 vdd3i! 17 19 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.54046e-13 AS=6.768e-13 PD=2.58169e-06 PS=3.78e-06 $X=620 $Y=2410 $dt=1
M19 17 RN vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.136e-13 AS=2.31854e-13 PD=2.4e-06 PS=1.31831e-06 $X=1460 $Y=2670 $dt=1
M20 23 19 vdd3i! vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=5.1875e-13 PD=6.7e-07 PS=2.99e-06 $X=3080 $Y=3400 $dt=1
M21 17 15 23 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=1.21617e-13 AS=5.25e-14 PD=9.13043e-07 PS=6.7e-07 $X=3630 $Y=3400 $dt=1
M22 22 9 17 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=1.2e-13 AS=2.77983e-13 PD=1.21e-06 PS=2.08696e-06 $X=4470 $Y=2860 $dt=1
M23 vdd3i! D 22 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=5.00229e-13 AS=1.2e-13 PD=2.34286e-06 PS=1.21e-06 $X=5020 $Y=2860 $dt=1
M24 15 C vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=4.94875e-13 AS=3.75171e-13 PD=3.04e-06 PS=1.75714e-06 $X=6060 $Y=2860 $dt=1
M25 vdd3i! 15 9 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.92547e-13 AS=3.528e-13 PD=1.8586e-06 PS=2.42e-06 $X=7720 $Y=2670 $dt=1
M26 21 19 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=1.25e-13 AS=5.45203e-13 PD=1.25e-06 PS=2.5814e-06 $X=8740 $Y=2820 $dt=1
M27 13 15 21 vdd3i! pe3i L=3e-07 W=1e-06 AD=2.96338e-13 AS=1.25e-13 PD=2.19718e-06 PS=1.25e-06 $X=9290 $Y=2820 $dt=1
M28 20 9 13 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=1.24462e-13 PD=6.7e-07 PS=9.22817e-07 $X=10150 $Y=3235 $dt=1
M29 vdd3i! 11 20 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=2.90656e-13 AS=5.25e-14 PD=1.25671e-06 PS=6.7e-07 $X=10700 $Y=3235 $dt=1
M30 vdd3i! RN 13 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=4.98268e-13 AS=2.976e-13 PD=2.15435e-06 PS=2.4e-06 $X=11900 $Y=2410 $dt=1
M31 11 13 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=9.75775e-13 PD=3.78e-06 PS=4.21894e-06 $X=12740 $Y=2410 $dt=1
M32 Q 13 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=1.1618e-12 PD=1.95e-06 PS=4.88e-06 $X=14480 $Y=2410 $dt=1
M33 vdd3i! 13 Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=3.807e-13 PD=1.95e-06 PS=1.95e-06 $X=15320 $Y=2410 $dt=1
M34 Q 13 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=3.807e-13 PD=1.95e-06 PS=1.95e-06 $X=16160 $Y=2410 $dt=1
M35 vdd3i! 13 Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=3.807e-13 PD=3.78e-06 PS=1.95e-06 $X=17000 $Y=2410 $dt=1
.ends DFRRQJI3VX4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX1 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=4
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.44533e-13 AS=2.016e-13 PD=1.44667e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=6.6e-07 AD=2.88e-13 AS=3.84267e-13 PD=2.28e-06 PS=2.27333e-06 $X=1590 $Y=890 $dt=0
M2 vdd3i! A 6 vdd3i! pe3i L=3e-07 W=9e-07 AD=4.7931e-13 AS=4.32e-13 PD=1.95649e-06 PS=2.76e-06 $X=620 $Y=2410 $dt=1
M3 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=5.712e-13 AS=7.7739e-13 PD=3.70971e-06 PS=3.17322e-06 $X=1640 $Y=2410 $dt=1
.ends BUJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO3I2JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO3I2JI3VX1 vdd3i! gnd3i! AN BN C Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 8 AN 9 gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=6e-14 AS=2.304e-13 PD=7.3e-07 PS=1.92e-06 $X=620 $Y=1070 $dt=0
M1 gnd3i! BN 8 gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=1.98937e-13 AS=6e-14 PD=1.31617e-06 PS=7.3e-07 $X=1220 $Y=1070 $dt=0
M2 Q C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.68863e-13 PD=1.43e-06 PS=2.4404e-06 $X=2060 $Y=660 $dt=0
M3 gnd3i! 9 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.329e-13 AS=2.403e-13 PD=2.77e-06 PS=1.43e-06 $X=2950 $Y=660 $dt=0
M4 9 AN vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=5.71409e-13 PD=1.24e-06 PS=2.5758e-06 $X=560 $Y=2590 $dt=1
M5 vdd3i! BN 9 vdd3i! pe3i L=3e-07 W=7e-07 AD=5.71409e-13 AS=1.89e-13 PD=2.5758e-06 PS=1.24e-06 $X=1400 $Y=2590 $dt=1
M6 10 C vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=1.15098e-12 PD=1.66e-06 PS=5.1884e-06 $X=2330 $Y=2410 $dt=1
M7 Q 9 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=8.46e-13 AS=1.7625e-13 PD=4.02e-06 PS=1.66e-06 $X=2880 $Y=2410 $dt=1
.ends NO3I2JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: FAJI3VX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt FAJI3VX1 vdd3i! gnd3i! S CI B A CO
*.DEVICECLIMB
** N=20 EP=7 FDC=28
M0 gnd3i! 12 S gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.361e-13 AS=4.272e-13 PD=2.76e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 15 CI 12 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=7.375e-14 AS=2.832e-13 PD=8.4e-07 PS=2.14e-06 $X=2220 $Y=960 $dt=0
M2 14 B 15 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=7.375e-14 AS=7.375e-14 PD=8.4e-07 PS=8.4e-07 $X=2820 $Y=960 $dt=0
M3 gnd3i! A 14 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=2.34033e-13 AS=7.375e-14 PD=1.52158e-06 PS=8.4e-07 $X=3420 $Y=960 $dt=0
M4 13 CI gnd3i! gnd3i! ne3i L=3.5e-07 W=5.5e-07 AD=1.485e-13 AS=2.18167e-13 PD=1.09e-06 PS=1.41842e-06 $X=4350 $Y=660 $dt=0
M5 gnd3i! A 13 gnd3i! ne3i L=3.5e-07 W=5.5e-07 AD=2.5017e-13 AS=1.485e-13 PD=1.58058e-06 PS=1.09e-06 $X=5240 $Y=660 $dt=0
M6 13 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=1.296e-13 AS=2.1833e-13 PD=1.02e-06 PS=1.37942e-06 $X=6220 $Y=960 $dt=0
M7 12 10 13 gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=2.304e-13 AS=1.296e-13 PD=1.92e-06 PS=1.02e-06 $X=7110 $Y=960 $dt=0
M8 gnd3i! 10 CO gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=3.345e-13 AS=2.832e-13 PD=1.73e-06 PS=2.14e-06 $X=8700 $Y=960 $dt=0
M9 11 A gnd3i! gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=7.375e-14 AS=3.345e-13 PD=8.4e-07 PS=1.73e-06 $X=9830 $Y=960 $dt=0
M10 10 B 11 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=1.593e-13 AS=7.375e-14 PD=1.13e-06 PS=8.4e-07 $X=10430 $Y=960 $dt=0
M11 9 CI 10 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=1.593e-13 AS=1.593e-13 PD=1.13e-06 PS=1.13e-06 $X=11320 $Y=960 $dt=0
M12 gnd3i! B 9 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=4.382e-13 AS=1.593e-13 PD=1.95e-06 PS=1.13e-06 $X=12210 $Y=960 $dt=0
M13 9 A gnd3i! gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=3.068e-13 AS=4.382e-13 PD=2.22e-06 PS=1.95e-06 $X=13550 $Y=960 $dt=0
M14 vdd3i! 12 S vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.6395e-13 AS=7.1205e-13 PD=4.52213e-06 PS=3.83e-06 $X=645 $Y=2410 $dt=1
M15 vdd3i! CI 17 vdd3i! pe3i L=3e-07 W=1.03e-06 AD=4.8155e-13 AS=4.79437e-13 PD=2.35e-06 PS=3.03778e-06 $X=2125 $Y=2490 $dt=1
M16 17 B vdd3i! vdd3i! pe3i L=3e-07 W=1.03e-06 AD=3.0385e-13 AS=4.8155e-13 PD=1.62e-06 PS=2.35e-06 $X=3095 $Y=2490 $dt=1
M17 vdd3i! A 17 vdd3i! pe3i L=3e-07 W=1.03e-06 AD=4.1015e-13 AS=3.0385e-13 PD=2.01e-06 PS=1.62e-06 $X=3985 $Y=2490 $dt=1
M18 20 A vdd3i! vdd3i! pe3i L=3e-07 W=1.03e-06 AD=1.545e-13 AS=4.1015e-13 PD=1.33e-06 PS=2.01e-06 $X=4955 $Y=2490 $dt=1
M19 19 B 20 vdd3i! pe3i L=3e-07 W=1.03e-06 AD=1.545e-13 AS=1.545e-13 PD=1.33e-06 PS=1.33e-06 $X=5555 $Y=2490 $dt=1
M20 12 CI 19 vdd3i! pe3i L=3e-07 W=1.03e-06 AD=3.0385e-13 AS=1.545e-13 PD=1.62e-06 PS=1.33e-06 $X=6155 $Y=2490 $dt=1
M21 17 10 12 vdd3i! pe3i L=3e-07 W=1.03e-06 AD=6.9155e-13 AS=3.0385e-13 PD=3.77e-06 PS=1.62e-06 $X=7045 $Y=2490 $dt=1
M22 vdd3i! 10 CO vdd3i! pe3i L=3e-07 W=1.11e-06 AD=4.54624e-13 AS=5.6055e-13 PD=2.27286e-06 PS=3.23e-06 $X=8675 $Y=2410 $dt=1
M23 16 A vdd3i! vdd3i! pe3i L=3e-07 W=9.9e-07 AD=2.9205e-13 AS=4.05476e-13 PD=1.58e-06 PS=2.02714e-06 $X=9645 $Y=2530 $dt=1
M24 vdd3i! B 16 vdd3i! pe3i L=3e-07 W=9.9e-07 AD=5.763e-13 AS=2.9205e-13 PD=3.59e-06 PS=1.58e-06 $X=10535 $Y=2530 $dt=1
M25 10 CI 16 vdd3i! pe3i L=3e-07 W=1e-06 AD=2.95e-13 AS=4.65e-13 PD=1.59e-06 PS=3.01e-06 $X=12085 $Y=2520 $dt=1
M26 18 B 10 vdd3i! pe3i L=3e-07 W=1e-06 AD=1.5e-13 AS=2.95e-13 PD=1.3e-06 PS=1.59e-06 $X=12975 $Y=2520 $dt=1
M27 vdd3i! A 18 vdd3i! pe3i L=3e-07 W=1e-06 AD=8.18e-13 AS=1.5e-13 PD=4.39e-06 PS=1.3e-06 $X=13575 $Y=2520 $dt=1
.ends FAJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OR2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OR2JI3VX0 vdd3i! gnd3i! A B Q
*.DEVICECLIMB
** N=8 EP=5 FDC=6
M0 7 A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.75467e-13 PD=9.6e-07 PS=2.95333e-06 $X=530 $Y=1130 $dt=0
M1 gnd3i! B 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.75467e-13 AS=1.134e-13 PD=2.95333e-06 PS=9.6e-07 $X=1420 $Y=1130 $dt=0
M2 Q 7 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=5.75467e-13 PD=1.8e-06 PS=2.95333e-06 $X=2390 $Y=1130 $dt=0
M3 8 A 7 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=4.08e-13 PD=1.1e-06 PS=2.66e-06 $X=620 $Y=2410 $dt=1
M4 vdd3i! B 8 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=8.28174e-13 AS=1.0625e-13 PD=2.99419e-06 PS=1.1e-06 $X=1170 $Y=2410 $dt=1
M5 Q 7 vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=3.36e-13 AS=6.82026e-13 PD=2.36e-06 PS=2.46581e-06 $X=2440 $Y=2410 $dt=1
.ends OR2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA3I1JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA3I1JI3VX1 vdd3i! gnd3i! AN Q B C
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 gnd3i! AN 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.40779e-13 AS=2.016e-13 PD=1.24397e-06 PS=1.8e-06 $X=620 $Y=660 $dt=0
M1 9 10 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.26825e-13 AS=5.10221e-13 PD=1.175e-06 PS=2.63603e-06 $X=1670 $Y=660 $dt=0
M2 8 B 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.31275e-13 AS=1.26825e-13 PD=1.185e-06 PS=1.175e-06 $X=2305 $Y=660 $dt=0
M3 Q C 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=1.31275e-13 PD=2.74e-06 PS=1.185e-06 $X=2950 $Y=660 $dt=0
M4 vdd3i! AN 10 vdd3i! pe3i L=3e-07 W=7e-07 AD=4.82246e-13 AS=3.36e-13 PD=2.26063e-06 PS=2.36e-06 $X=620 $Y=2410 $dt=1
M5 vdd3i! 10 Q vdd3i! pe3i L=3.00059e-07 W=1.00314e-06 AD=6.91085e-13 AS=2.195e-13 PD=3.2396e-06 PS=1.46314e-06 $X=1430 $Y=2410 $dt=1
M6 Q B vdd3i! vdd3i! pe3i L=3.00059e-07 W=1.00314e-06 AD=2.195e-13 AS=6.91085e-13 PD=1.46314e-06 PS=3.2396e-06 $X=2270 $Y=2410 $dt=1
M7 Q C vdd3i! vdd3i! pe3i L=3.00059e-07 W=1.00314e-06 AD=4.232e-13 AS=6.91085e-13 PD=2.85314e-06 PS=3.2396e-06 $X=3000 $Y=2410 $dt=1
.ends NA3I1JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DLY2JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DLY2JI3VX1 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=12 EP=4 FDC=12
M0 gnd3i! A 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.577e-13 AS=2.016e-13 PD=1.79e-06 PS=1.8e-06 $X=620 $Y=660 $dt=0
M1 8 10 gnd3i! gnd3i! ne3i L=8e-07 W=4.2e-07 AD=2.548e-13 AS=3.577e-13 PD=1.7e-06 PS=1.79e-06 $X=1990 $Y=660 $dt=0
M2 8 10 9 gnd3i! ne3i L=8e-07 W=4.2e-07 AD=2.548e-13 AS=2.016e-13 PD=1.7e-06 PS=1.8e-06 $X=1990 $Y=1360 $dt=0
M3 gnd3i! 9 7 gnd3i! ne3i L=1e-06 W=4.2e-07 AD=3.42444e-13 AS=2.1e-13 PD=1.66718e-06 PS=1.62e-06 $X=3950 $Y=660 $dt=0
M4 6 9 7 gnd3i! ne3i L=1e-06 W=4.2e-07 AD=2.10588e-13 AS=2.1e-13 PD=1.81778e-06 PS=1.62e-06 $X=3950 $Y=1360 $dt=0
M5 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=7.25656e-13 PD=2.74e-06 PS=3.53282e-06 $X=6310 $Y=660 $dt=0
M6 vdd3i! A 10 vdd3i! pe3i L=3e-07 W=7e-07 AD=5.42937e-13 AS=3.535e-13 PD=2.69375e-06 PS=2.41e-06 $X=645 $Y=3120 $dt=1
M7 12 10 9 vdd3i! pe3i L=7.4e-07 W=4.2e-07 AD=2.8095e-13 AS=2.0035e-13 PD=1.785e-06 PS=1.77071e-06 $X=2050 $Y=2640 $dt=1
M8 12 10 vdd3i! vdd3i! pe3i L=7.4e-07 W=4.2e-07 AD=2.8095e-13 AS=3.25762e-13 PD=1.785e-06 PS=1.61625e-06 $X=2050 $Y=3400 $dt=1
M9 6 9 11 vdd3i! pe3i L=1e-06 W=4.2e-07 AD=2.856e-13 AS=2.479e-13 PD=2.2e-06 PS=1.715e-06 $X=4030 $Y=2660 $dt=1
M10 vdd3i! 9 11 vdd3i! pe3i L=1e-06 W=4.2e-07 AD=2.62018e-13 AS=2.479e-13 PD=1.40689e-06 PS=1.715e-06 $X=4030 $Y=3400 $dt=1
M11 Q 6 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.1205e-13 AS=8.79632e-13 PD=3.83e-06 PS=4.72311e-06 $X=6335 $Y=2410 $dt=1
.ends DLY2JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA3JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA3JI3VX0 vdd3i! gnd3i! C Q B A
*.DEVICECLIMB
** N=9 EP=6 FDC=6
M0 9 C gnd3i! gnd3i! ne3i L=3.5e-07 W=7e-07 AD=8.75e-14 AS=5.605e-13 PD=9.5e-07 PS=3.52e-06 $X=630 $Y=850 $dt=0
M1 8 B 9 gnd3i! ne3i L=3.5e-07 W=7e-07 AD=8.75e-14 AS=8.75e-14 PD=9.5e-07 PS=9.5e-07 $X=1230 $Y=850 $dt=0
M2 Q A 8 gnd3i! ne3i L=3.5e-07 W=7e-07 AD=3.36e-13 AS=8.75e-14 PD=2.36e-06 PS=9.5e-07 $X=1830 $Y=850 $dt=0
M3 Q C vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=5.76467e-13 PD=1.24e-06 PS=3.21333e-06 $X=470 $Y=2580 $dt=1
M4 vdd3i! B Q vdd3i! pe3i L=3e-07 W=7e-07 AD=5.76467e-13 AS=1.89e-13 PD=3.21333e-06 PS=1.24e-06 $X=1310 $Y=2580 $dt=1
M5 Q A vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=4.708e-13 AS=5.76467e-13 PD=3.92e-06 PS=3.21333e-06 $X=2040 $Y=2470 $dt=1
.ends NA3JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ON21JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ON21JI3VX1 vdd3i! gnd3i! B A Q C
*.DEVICECLIMB
** N=9 EP=6 FDC=6
M0 gnd3i! B 8 gnd3i! ne3i L=3.4958e-07 W=8.92071e-07 AD=2.40125e-13 AS=4.24712e-13 PD=1.43207e-06 PS=2.73707e-06 $X=615 $Y=660 $dt=0
M1 8 A gnd3i! gnd3i! ne3i L=3.4958e-07 W=8.92071e-07 AD=2.37987e-13 AS=2.40125e-13 PD=1.42707e-06 PS=1.43207e-06 $X=1505 $Y=660 $dt=0
M2 Q C 8 gnd3i! ne3i L=3.4958e-07 W=8.92071e-07 AD=4.24712e-13 AS=2.37987e-13 PD=2.73707e-06 PS=1.42707e-06 $X=2395 $Y=660 $dt=0
M3 9 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=9.418e-13 PD=1.66e-06 PS=4.63e-06 $X=695 $Y=2410 $dt=1
M4 Q A 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.75706e-13 AS=1.7625e-13 PD=2.44322e-06 PS=1.66e-06 $X=1245 $Y=2410 $dt=1
M5 vdd3i! C Q vdd3i! pe3i L=3e-07 W=9.85e-07 AD=1.1721e-12 AS=3.32319e-13 PD=4.94e-06 PS=1.70678e-06 $X=2210 $Y=2410 $dt=1
.ends ON21JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OA21JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OA21JI3VX1 vdd3i! gnd3i! C A B Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 8 C 9 gnd3i! ne3i L=3.5e-07 W=5.4e-07 AD=3.313e-13 AS=2.97e-13 PD=1.95333e-06 PS=2.18e-06 $X=690 $Y=660 $dt=0
M1 8 A gnd3i! gnd3i! ne3i L=3.5e-07 W=5.4e-07 AD=3.313e-13 AS=2.592e-13 PD=1.95333e-06 PS=2.04e-06 $X=1620 $Y=1480 $dt=0
M2 gnd3i! B 8 gnd3i! ne3i L=3.5e-07 W=5.4e-07 AD=2.92808e-13 AS=3.313e-13 PD=1.47273e-06 PS=1.95333e-06 $X=2450 $Y=1010 $dt=0
M3 Q 9 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=4.82592e-13 PD=2.74e-06 PS=2.42727e-06 $X=3510 $Y=660 $dt=0
M4 9 C vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=2.295e-13 AS=1.03315e-12 PD=1.39e-06 PS=4.25e-06 $X=975 $Y=2880 $dt=1
M5 10 A 9 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=2.295e-13 PD=1.1e-06 PS=1.39e-06 $X=1815 $Y=2880 $dt=1
M6 vdd3i! B 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.77448e-13 AS=1.0625e-13 PD=1.94425e-06 PS=1.1e-06 $X=2365 $Y=2880 $dt=1
M7 Q 9 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=7.92002e-13 PD=3.78e-06 PS=3.22516e-06 $X=3560 $Y=2410 $dt=1
.ends OA21JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX3                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX3 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=7
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=5.23e-13 AS=4.272e-13 PD=2.14e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.5365e-13 AS=5.23e-13 PD=1.46e-06 PS=2.14e-06 $X=1870 $Y=660 $dt=0
M2 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=7.586e-13 AS=2.5365e-13 PD=3.76e-06 PS=1.46e-06 $X=2790 $Y=660 $dt=0
M3 vdd3i! A 6 vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=6.11825e-13 AS=5.712e-13 PD=2.51971e-06 PS=3.70971e-06 $X=620 $Y=2410 $dt=1
M4 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=6.11825e-13 PD=1.87971e-06 PS=2.51971e-06 $X=1510 $Y=2410 $dt=1
M5 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=3.3675e-13 AS=2.751e-13 PD=1.92971e-06 PS=1.87971e-06 $X=2350 $Y=2410 $dt=1
M6 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=5.712e-13 AS=3.3675e-13 PD=3.70971e-06 PS=1.92971e-06 $X=3000 $Y=2410 $dt=1
.ends BUJI3VX3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AN211JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AN211JI3VX1 vdd3i! gnd3i! B A Q C D
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 9 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=6.47e-13 PD=1.14e-06 PS=3.58e-06 $X=690 $Y=660 $dt=0
M1 Q A 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.9785e-13 AS=1.1125e-13 PD=1.71704e-06 PS=1.14e-06 $X=1290 $Y=660 $dt=0
M2 gnd3i! C Q gnd3i! ne3i L=3.5e-07 W=6.65e-07 AD=5.036e-13 AS=2.2255e-13 PD=2.145e-06 PS=1.28296e-06 $X=2250 $Y=885 $dt=0
M3 Q D gnd3i! gnd3i! ne3i L=3.5e-07 W=6.65e-07 AD=3.22525e-13 AS=5.036e-13 PD=2.3e-06 PS=2.145e-06 $X=3505 $Y=885 $dt=0
M4 vdd3i! B 11 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.5825e-13 AS=6.768e-13 PD=2.06e-06 PS=3.78e-06 $X=620 $Y=2410 $dt=1
M5 11 A vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=4.5825e-13 PD=2e-06 PS=2.06e-06 $X=1570 $Y=2410 $dt=1
M6 10 C 11 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.115e-13 AS=4.1595e-13 PD=1.71e-06 PS=2e-06 $X=2460 $Y=2410 $dt=1
M7 Q D 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=2.115e-13 PD=3.78e-06 PS=1.71e-06 $X=3060 $Y=2410 $dt=1
.ends AN211JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX16                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX16 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=39
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=4.272e-13 PD=1.43e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=1510 $Y=660 $dt=0
M2 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=2400 $Y=660 $dt=0
M3 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=3290 $Y=660 $dt=0
M4 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=4180 $Y=660 $dt=0
M5 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.4475e-13 AS=2.403e-13 PD=1.44e-06 PS=1.43e-06 $X=5070 $Y=660 $dt=0
M6 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.63267e-13 AS=2.4475e-13 PD=1.95905e-06 PS=1.44e-06 $X=5970 $Y=660 $dt=0
M7 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.26533e-13 PD=1.34e-06 PS=1.76095e-06 $X=6940 $Y=750 $dt=0
M8 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=7830 $Y=750 $dt=0
M9 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=8800 $Y=750 $dt=0
M10 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=9690 $Y=750 $dt=0
M11 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=10660 $Y=750 $dt=0
M12 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=11550 $Y=750 $dt=0
M13 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=12520 $Y=750 $dt=0
M14 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=13410 $Y=750 $dt=0
M15 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=14380 $Y=750 $dt=0
M16 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.84e-13 AS=2.16e-13 PD=2.56e-06 PS=1.34e-06 $X=15270 $Y=750 $dt=0
M17 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=5.79287e-13 PD=1.86506e-06 PS=3.69506e-06 $X=475 $Y=2410 $dt=1
M18 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1315 $Y=2410 $dt=1
M19 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1865 $Y=2410 $dt=1
M20 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=2705 $Y=2410 $dt=1
M21 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=3255 $Y=2410 $dt=1
M22 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=4095 $Y=2410 $dt=1
M23 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=4645 $Y=2410 $dt=1
M24 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=5485 $Y=2410 $dt=1
M25 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=6035 $Y=2410 $dt=1
M26 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=6875 $Y=2410 $dt=1
M27 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=7425 $Y=2410 $dt=1
M28 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=8265 $Y=2410 $dt=1
M29 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=8815 $Y=2410 $dt=1
M30 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=9655 $Y=2410 $dt=1
M31 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=10205 $Y=2410 $dt=1
M32 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=11045 $Y=2410 $dt=1
M33 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=11595 $Y=2410 $dt=1
M34 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=12435 $Y=2410 $dt=1
M35 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=12985 $Y=2410 $dt=1
M36 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=13825 $Y=2410 $dt=1
M37 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=14375 $Y=2410 $dt=1
M38 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=1.15229e-12 AS=2.54913e-13 PD=4.89506e-06 PS=1.86506e-06 $X=15215 $Y=2410 $dt=1
.ends BUJI3VX16

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX0                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX0 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=4
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.923e-13 AS=2.016e-13 PD=2.005e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=3.923e-13 PD=1.8e-06 PS=2.005e-06 $X=1735 $Y=1130 $dt=0
M2 vdd3i! A 6 vdd3i! pe3i L=3e-07 W=9e-07 AD=5.7805e-13 AS=4.32e-13 PD=2.33911e-06 PS=2.76e-06 $X=620 $Y=2410 $dt=1
M3 Q 6 vdd3i! vdd3i! pe3i L=3e-07 W=1.12e-06 AD=5.376e-13 AS=7.1935e-13 PD=3.2e-06 PS=2.91089e-06 $X=1785 $Y=2410 $dt=1
.ends BUJI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA2I1JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA2I1JI3VX1 vdd3i! gnd3i! AN Q B
*.DEVICECLIMB
** N=8 EP=5 FDC=6
M0 gnd3i! AN 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.44754e-13 AS=2.016e-13 PD=1.25038e-06 PS=1.8e-06 $X=620 $Y=660 $dt=0
M1 7 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=5.18646e-13 PD=1.14e-06 PS=2.64962e-06 $X=1680 $Y=660 $dt=0
M2 Q B 7 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=1.1125e-13 PD=2.74e-06 PS=1.14e-06 $X=2280 $Y=660 $dt=0
M3 vdd3i! AN 8 vdd3i! pe3i L=3e-07 W=7e-07 AD=6.84341e-13 AS=3.36e-13 PD=3.08e-06 PS=2.36e-06 $X=620 $Y=2410 $dt=1
M4 Q 8 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.7e-13 AS=9.7763e-13 PD=1.54e-06 PS=4.4e-06 $X=1510 $Y=2410 $dt=1
M5 vdd3i! B Q vdd3i! pe3i L=3e-07 W=1e-06 AD=9.7763e-13 AS=2.7e-13 PD=4.4e-06 PS=1.54e-06 $X=2350 $Y=2410 $dt=1
.ends NA2I1JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DLY1JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DLY1JI3VX1 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=8 EP=4 FDC=8
M0 gnd3i! A 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.591e-13 AS=2.016e-13 PD=2.13e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 6 8 gnd3i! gnd3i! ne3i L=8e-07 W=4.2e-07 AD=2.415e-13 AS=3.591e-13 PD=1.99e-06 PS=2.13e-06 $X=1590 $Y=1400 $dt=0
M2 gnd3i! 6 7 gnd3i! ne3i L=1e-06 W=4.2e-07 AD=2.6662e-13 AS=2.016e-13 PD=1.28565e-06 PS=1.8e-06 $X=2860 $Y=660 $dt=0
M3 Q 7 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.3165e-13 AS=5.6498e-13 PD=2.75e-06 PS=2.72435e-06 $X=4625 $Y=660 $dt=0
M4 vdd3i! A 8 vdd3i! pe3i L=3e-07 W=6.7e-07 AD=4.61962e-13 AS=3.3835e-13 PD=2.62468e-06 PS=2.35e-06 $X=645 $Y=2680 $dt=1
M5 6 8 vdd3i! vdd3i! pe3i L=1e-06 W=4.2e-07 AD=2.00088e-13 AS=2.89588e-13 PD=1.76778e-06 PS=1.64532e-06 $X=1590 $Y=2680 $dt=1
M6 vdd3i! 6 7 vdd3i! pe3i L=7.5e-07 W=4.2e-07 AD=2.78313e-13 AS=2.00088e-13 PD=1.17049e-06 PS=1.76778e-06 $X=3110 $Y=3400 $dt=1
M7 Q 7 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.191e-13 AS=9.34337e-13 PD=3.84e-06 PS=3.92951e-06 $X=4650 $Y=2410 $dt=1
.ends DLY1JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OR4JI3VX1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OR4JI3VX1 vdd3i! gnd3i! C D Q B A
*.DEVICECLIMB
** N=13 EP=7 FDC=12
M0 11 C gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=4.12474e-13 PD=9.6e-07 PS=2.12185e-06 $X=510 $Y=1130 $dt=0
M1 gnd3i! D 11 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=4.12474e-13 AS=1.134e-13 PD=2.12185e-06 PS=9.6e-07 $X=1400 $Y=1130 $dt=0
M2 10 11 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=8.74052e-13 PD=1.14e-06 PS=4.4963e-06 $X=2330 $Y=660 $dt=0
M3 Q 9 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.56e-13 AS=1.1125e-13 PD=2.64627e-06 PS=1.14e-06 $X=2930 $Y=660 $dt=0
M4 9 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=7.908e-13 PD=9.6e-07 PS=4.27314e-06 $X=4410 $Y=1130 $dt=0
M5 gnd3i! A 9 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=7.908e-13 AS=1.134e-13 PD=4.27314e-06 PS=9.6e-07 $X=5300 $Y=1130 $dt=0
M6 13 C 11 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=4.08e-13 PD=1.1e-06 PS=2.66e-06 $X=620 $Y=2410 $dt=1
M7 vdd3i! D 13 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=6.21177e-13 AS=1.0625e-13 PD=2.08363e-06 PS=1.1e-06 $X=1170 $Y=2410 $dt=1
M8 Q 11 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=1.03042e-12 PD=1.95e-06 PS=3.45637e-06 $X=2480 $Y=2410 $dt=1
M9 vdd3i! 9 Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.09631e-12 AS=3.807e-13 PD=3.53124e-06 PS=1.95e-06 $X=3320 $Y=2410 $dt=1
M10 12 B vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=6.60894e-13 PD=1.1e-06 PS=2.12876e-06 $X=4690 $Y=2410 $dt=1
M11 9 A 12 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.08e-13 AS=1.0625e-13 PD=2.66e-06 PS=1.1e-06 $X=5240 $Y=2410 $dt=1
.ends OR4JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DFRRQJI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DFRRQJI3VX1 vdd3i! gnd3i! RN D C Q
*.DEVICECLIMB
** N=23 EP=6 FDC=30
M0 gnd3i! 17 19 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.39017e-13 AS=2.016e-13 PD=9.16947e-07 PS=1.8e-06 $X=620 $Y=660 $dt=0
M1 10 RN gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.28952e-13 AS=2.94583e-13 PD=2.36956e-06 PS=1.94305e-06 $X=1510 $Y=660 $dt=0
M2 18 19 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.55236e-13 PD=6.7e-07 PS=1.11822e-06 $X=2340 $Y=1390 $dt=0
M3 17 9 18 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=2940 $Y=1390 $dt=0
M4 16 15 17 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=3830 $Y=1390 $dt=0
M5 10 D 16 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.835e-13 AS=5.25e-14 PD=2.19e-06 PS=6.7e-07 $X=4430 $Y=1390 $dt=0
M6 gnd3i! C 15 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.659e-13 AS=2.016e-13 PD=1.21e-06 PS=1.8e-06 $X=6060 $Y=1390 $dt=0
M7 9 15 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.95e-13 AS=1.659e-13 PD=2.23e-06 PS=1.21e-06 $X=7045 $Y=1390 $dt=0
M8 14 19 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=8695 $Y=1020 $dt=0
M9 13 9 14 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=9295 $Y=1020 $dt=0
M10 12 15 13 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=10185 $Y=1020 $dt=0
M11 8 11 12 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.55817e-13 AS=5.25e-14 PD=9.68244e-07 PS=6.7e-07 $X=10785 $Y=1020 $dt=0
M12 gnd3i! RN 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=6.52289e-13 AS=3.30183e-13 PD=3.3375e-06 PS=2.05176e-06 $X=11755 $Y=660 $dt=0
M13 11 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=3.07822e-13 PD=1.8e-06 PS=1.575e-06 $X=12560 $Y=1130 $dt=0
M14 Q 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=6.52289e-13 PD=2.74e-06 PS=3.3375e-06 $X=14150 $Y=660 $dt=0
M15 vdd3i! 17 19 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=1.944e-13 AS=3.456e-13 PD=1.26e-06 PS=2.4e-06 $X=620 $Y=2670 $dt=1
M16 17 RN vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.136e-13 AS=1.944e-13 PD=2.4e-06 PS=1.26e-06 $X=1460 $Y=2670 $dt=1
M17 23 19 vdd3i! vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=5.1875e-13 PD=6.7e-07 PS=2.99e-06 $X=3080 $Y=3400 $dt=1
M18 17 15 23 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=1.21617e-13 AS=5.25e-14 PD=9.13043e-07 PS=6.7e-07 $X=3630 $Y=3400 $dt=1
M19 22 9 17 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=1.2e-13 AS=2.77983e-13 PD=1.21e-06 PS=2.08696e-06 $X=4470 $Y=2860 $dt=1
M20 vdd3i! D 22 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=5.00229e-13 AS=1.2e-13 PD=2.34286e-06 PS=1.21e-06 $X=5020 $Y=2860 $dt=1
M21 15 C vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=4.94875e-13 AS=3.75171e-13 PD=3.04e-06 PS=1.75714e-06 $X=6060 $Y=2860 $dt=1
M22 vdd3i! 15 9 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.92547e-13 AS=3.528e-13 PD=1.8586e-06 PS=2.42e-06 $X=7720 $Y=2670 $dt=1
M23 21 19 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=1.25e-13 AS=5.45203e-13 PD=1.25e-06 PS=2.5814e-06 $X=8740 $Y=2820 $dt=1
M24 13 15 21 vdd3i! pe3i L=3e-07 W=1e-06 AD=2.96338e-13 AS=1.25e-13 PD=2.19718e-06 PS=1.25e-06 $X=9290 $Y=2820 $dt=1
M25 20 9 13 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=1.24462e-13 PD=6.7e-07 PS=9.22817e-07 $X=10150 $Y=3235 $dt=1
M26 vdd3i! 11 20 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=4.10996e-13 AS=5.25e-14 PD=1.64789e-06 PS=6.7e-07 $X=10700 $Y=3235 $dt=1
M27 vdd3i! RN 13 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=7.04565e-13 AS=2.976e-13 PD=2.82495e-06 PS=2.4e-06 $X=11900 $Y=2410 $dt=1
M28 11 13 vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.456e-13 AS=7.04565e-13 PD=2.4e-06 PS=2.82495e-06 $X=12740 $Y=2410 $dt=1
M29 Q 13 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=1.37977e-12 PD=3.78e-06 PS=5.5322e-06 $X=14200 $Y=2410 $dt=1
.ends DFRRQJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INJI3VX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INJI3VX1 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=5 EP=4 FDC=2
M0 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=6e-07 AD=2.88e-13 AS=6.428e-13 PD=2.16e-06 PS=3.62e-06 $X=710 $Y=950 $dt=0
M1 Q A vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=1.0562e-12 PD=3.78e-06 PS=4.76e-06 $X=760 $Y=2410 $dt=1
.ends INJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INJI3VX2                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INJI3VX2 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=5 EP=4 FDC=4
M0 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=1.296e-13 AS=4.408e-13 PD=1.02e-06 PS=3.52e-06 $X=500 $Y=1070 $dt=0
M1 gnd3i! A Q gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=4.408e-13 AS=1.296e-13 PD=3.52e-06 PS=1.02e-06 $X=1390 $Y=1070 $dt=0
M2 Q A vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=8.151e-13 PD=1.87971e-06 PS=4.50971e-06 $X=560 $Y=2410 $dt=1
M3 vdd3i! A Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=8.01e-13 AS=2.751e-13 PD=4.48971e-06 PS=1.87971e-06 $X=1400 $Y=2410 $dt=1
.ends INJI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX12                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX12 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=28
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=4.148e-13 AS=3.84e-13 PD=1.98e-06 PS=2.56e-06 $X=620 $Y=750 $dt=0
M1 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=4.148e-13 PD=1.34e-06 PS=1.98e-06 $X=1710 $Y=750 $dt=0
M2 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=2600 $Y=750 $dt=0
M3 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=3570 $Y=750 $dt=0
M4 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=4460 $Y=750 $dt=0
M5 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=5430 $Y=750 $dt=0
M6 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=6320 $Y=750 $dt=0
M7 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=7290 $Y=750 $dt=0
M8 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=8180 $Y=750 $dt=0
M9 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=9150 $Y=750 $dt=0
M10 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.194e-13 AS=2.16e-13 PD=1.36e-06 PS=1.34e-06 $X=10040 $Y=750 $dt=0
M11 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.84e-13 AS=2.194e-13 PD=2.56e-06 PS=1.36e-06 $X=10930 $Y=750 $dt=0
M12 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=5.79287e-13 PD=1.86506e-06 PS=3.69506e-06 $X=475 $Y=2410 $dt=1
M13 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1315 $Y=2410 $dt=1
M14 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1865 $Y=2410 $dt=1
M15 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=2705 $Y=2410 $dt=1
M16 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=3255 $Y=2410 $dt=1
M17 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=4095 $Y=2410 $dt=1
M18 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=4645 $Y=2410 $dt=1
M19 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=5485 $Y=2410 $dt=1
M20 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=6035 $Y=2410 $dt=1
M21 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=6875 $Y=2410 $dt=1
M22 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=7425 $Y=2410 $dt=1
M23 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=8265 $Y=2410 $dt=1
M24 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=8815 $Y=2410 $dt=1
M25 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=9655 $Y=2410 $dt=1
M26 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=10205 $Y=2410 $dt=1
M27 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=8.53088e-13 AS=2.54913e-13 PD=4.55506e-06 PS=1.86506e-06 $X=11045 $Y=2410 $dt=1
.ends BUJI3VX12

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ON22JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ON22JI3VX1 vdd3i! gnd3i! D C Q A B
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 gnd3i! D 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=4.272e-13 PD=1.86e-06 PS=2.74e-06 $X=720 $Y=660 $dt=0
M1 9 C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=1690 $Y=660 $dt=0
M2 Q A 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=2580 $Y=660 $dt=0
M3 9 B Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.666e-13 AS=2.403e-13 PD=2.84e-06 PS=1.43e-06 $X=3470 $Y=660 $dt=0
M4 11 D vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=8.802e-13 PD=1.66e-06 PS=4.56e-06 $X=1120 $Y=2410 $dt=1
M5 Q C 11 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=1.7625e-13 PD=1.95e-06 PS=1.66e-06 $X=1670 $Y=2410 $dt=1
M6 10 A Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=3.807e-13 PD=1.66e-06 PS=1.95e-06 $X=2510 $Y=2410 $dt=1
M7 vdd3i! B 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=8.802e-13 AS=1.7625e-13 PD=4.56e-06 PS=1.66e-06 $X=3060 $Y=2410 $dt=1
.ends ON22JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AN31JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AN31JI3VX1 vdd3i! gnd3i! A B C Q D
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 10 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.335e-13 AS=6.098e-13 PD=1.19e-06 PS=3.52e-06 $X=660 $Y=660 $dt=0
M1 9 B 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.35725e-13 AS=1.335e-13 PD=1.195e-06 PS=1.19e-06 $X=1310 $Y=660 $dt=0
M2 Q C 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.0257e-13 AS=1.35725e-13 PD=1.8043e-06 PS=1.195e-06 $X=1965 $Y=660 $dt=0
M3 gnd3i! D Q gnd3i! ne3i L=3.5e-07 W=5.75e-07 AD=5.783e-13 AS=1.9548e-13 PD=3.52e-06 PS=1.1657e-06 $X=2910 $Y=975 $dt=0
M4 11 A vdd3i! vdd3i! pe3i L=3.00061e-07 W=1.44471e-06 AD=3.0525e-13 AS=5.93475e-13 PD=1.86471e-06 PS=3.72971e-06 $X=525 $Y=2425 $dt=1
M5 vdd3i! B 11 vdd3i! pe3i L=3.00061e-07 W=1.44471e-06 AD=4.42387e-13 AS=3.0525e-13 PD=2.08971e-06 PS=1.86471e-06 $X=1365 $Y=2425 $dt=1
M6 11 C vdd3i! vdd3i! pe3i L=3.00061e-07 W=1.44471e-06 AD=2.6565e-13 AS=4.42387e-13 PD=1.86471e-06 PS=2.08971e-06 $X=2310 $Y=2425 $dt=1
M7 Q D 11 vdd3i! pe3i L=3.00061e-07 W=1.44471e-06 AD=7.2375e-13 AS=2.6565e-13 PD=3.85971e-06 PS=1.86471e-06 $X=2910 $Y=2425 $dt=1
.ends AN31JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO3JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO3JI3VX0 vdd3i! gnd3i! C Q B A
*.DEVICECLIMB
** N=9 EP=6 FDC=6
M0 Q C gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.75467e-13 PD=9.6e-07 PS=2.95333e-06 $X=615 $Y=1130 $dt=0
M1 gnd3i! B Q gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.75467e-13 AS=1.134e-13 PD=2.95333e-06 PS=9.6e-07 $X=1505 $Y=1130 $dt=0
M2 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=5.75467e-13 PD=1.8e-06 PS=2.95333e-06 $X=2390 $Y=1130 $dt=0
M3 9 C vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=1.55e-13 AS=1.3584e-12 PD=1.31e-06 PS=5.15e-06 $X=955 $Y=2410 $dt=1
M4 8 B 9 vdd3i! pe3i L=3e-07 W=1e-06 AD=1.55e-13 AS=1.55e-13 PD=1.31e-06 PS=1.31e-06 $X=1565 $Y=2410 $dt=1
M5 Q A 8 vdd3i! pe3i L=3e-07 W=1e-06 AD=4.8e-13 AS=1.55e-13 PD=2.96e-06 PS=1.31e-06 $X=2175 $Y=2410 $dt=1
.ends NO3JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OR4JI3VX2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OR4JI3VX2 vdd3i! gnd3i! C D Q B A
*.DEVICECLIMB
** N=14 EP=7 FDC=16
M0 10 C gnd3i! gnd3i! ne3i L=3.5e-07 W=7e-07 AD=1.9155e-13 AS=3.417e-13 PD=1.255e-06 PS=2.39e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! D 10 gnd3i! ne3i L=3.5e-07 W=7e-07 AD=2.07711e-13 AS=1.9155e-13 PD=1.27673e-06 PS=1.255e-06 $X=1510 $Y=660 $dt=0
M2 12 10 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=2.64089e-13 PD=1.14e-06 PS=1.62327e-06 $X=2420 $Y=660 $dt=0
M3 Q 9 12 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=1.1125e-13 PD=1.43e-06 PS=1.14e-06 $X=3020 $Y=660 $dt=0
M4 11 9 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.2015e-13 AS=2.403e-13 PD=1.16e-06 PS=1.43e-06 $X=3910 $Y=660 $dt=0
M5 gnd3i! 10 11 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.54126e-13 AS=1.2015e-13 PD=1.60088e-06 PS=1.16e-06 $X=4530 $Y=660 $dt=0
M6 9 B gnd3i! gnd3i! ne3i L=3.5e-07 W=7e-07 AD=1.9155e-13 AS=1.99874e-13 PD=1.255e-06 PS=1.25912e-06 $X=5420 $Y=660 $dt=0
M7 gnd3i! A 9 gnd3i! ne3i L=3.5e-07 W=7e-07 AD=3.417e-13 AS=1.9155e-13 PD=2.39e-06 PS=1.255e-06 $X=6310 $Y=660 $dt=0
M8 14 C 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=6.768e-13 PD=1.66e-06 PS=3.78e-06 $X=710 $Y=2410 $dt=1
M9 vdd3i! D 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=5.47043e-13 AS=1.7625e-13 PD=2.41704e-06 PS=1.66e-06 $X=1260 $Y=2410 $dt=1
M10 Q 10 vdd3i! vdd3i! pe3i L=2.99799e-07 W=1.41828e-06 AD=3.622e-13 AS=5.50257e-13 PD=1.93828e-06 PS=2.43124e-06 $X=2210 $Y=2410 $dt=1
M11 vdd3i! 9 Q vdd3i! pe3i L=2.99799e-07 W=1.41828e-06 AD=4.987e-13 AS=3.622e-13 PD=2.36828e-06 PS=1.93828e-06 $X=3050 $Y=2410 $dt=1
M12 Q 9 vdd3i! vdd3i! pe3i L=2.99799e-07 W=1.41828e-06 AD=3.622e-13 AS=4.987e-13 PD=1.93828e-06 PS=2.36828e-06 $X=3930 $Y=2410 $dt=1
M13 vdd3i! 10 Q vdd3i! pe3i L=2.99799e-07 W=1.41828e-06 AD=5.8556e-13 AS=3.622e-13 PD=2.47136e-06 PS=1.93828e-06 $X=4770 $Y=2410 $dt=1
M14 13 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=5.8214e-13 PD=1.66e-06 PS=2.45692e-06 $X=5760 $Y=2410 $dt=1
M15 9 A 13 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=1.7625e-13 PD=3.78e-06 PS=1.66e-06 $X=6310 $Y=2410 $dt=1
.ends OR4JI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: HAJI3VX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt HAJI3VX1 vdd3i! gnd3i! S B A CO
*.DEVICECLIMB
** N=12 EP=6 FDC=14
M0 gnd3i! 8 S gnd3i! ne3i L=3.49889e-07 W=8.98284e-07 AD=4.998e-13 AS=4.174e-13 PD=3.41456e-06 PS=2.72828e-06 $X=600 $Y=660 $dt=0
M1 gnd3i! A 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.52e-13 PD=1.43e-06 PS=2.74e-06 $X=2070 $Y=660 $dt=0
M2 9 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.70969e-13 AS=2.403e-13 PD=1.71986e-06 PS=1.43e-06 $X=2960 $Y=660 $dt=0
M3 8 10 9 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=3.632e-13 AS=1.79631e-13 PD=2.84284e-06 PS=1.14014e-06 $X=3850 $Y=960 $dt=0
M4 gnd3i! 10 CO gnd3i! ne3i L=3.5e-07 W=5.5e-07 AD=1.56292e-13 AS=2.4195e-13 PD=1.09236e-06 PS=2.03071e-06 $X=5380 $Y=1000 $dt=0
M5 11 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=2.52908e-13 PD=1.14e-06 PS=1.76764e-06 $X=6270 $Y=660 $dt=0
M6 10 A 11 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=1.1125e-13 PD=2.74e-06 PS=1.14e-06 $X=6870 $Y=660 $dt=0
M7 vdd3i! 8 S vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.07833e-13 AS=7.1205e-13 PD=2.97939e-06 PS=3.83e-06 $X=645 $Y=2410 $dt=1
M8 12 A vdd3i! vdd3i! pe3i L=3e-07 W=8.9e-07 AD=1.335e-13 AS=3.83667e-13 PD=1.19e-06 PS=1.88061e-06 $X=1615 $Y=2630 $dt=1
M9 8 B 12 vdd3i! pe3i L=3e-07 W=8.9e-07 AD=4.9565e-13 AS=1.335e-13 PD=2.12e-06 PS=1.19e-06 $X=2215 $Y=2630 $dt=1
M10 vdd3i! 10 8 vdd3i! pe3i L=3e-07 W=8.9e-07 AD=4.8925e-13 AS=4.9565e-13 PD=3.49e-06 PS=2.12e-06 $X=3525 $Y=2630 $dt=1
M11 vdd3i! 10 CO vdd3i! pe3i L=3e-07 W=1.11e-06 AD=4.3695e-13 AS=4.7415e-13 PD=2.09e-06 PS=3.23e-06 $X=4995 $Y=2410 $dt=1
M12 10 B vdd3i! vdd3i! pe3i L=3e-07 W=1.11e-06 AD=3.2745e-13 AS=4.3695e-13 PD=1.7e-06 PS=2.09e-06 $X=5965 $Y=2410 $dt=1
M13 vdd3i! A 10 vdd3i! pe3i L=3e-07 W=1.11e-06 AD=8.7795e-13 AS=3.2745e-13 PD=4.61e-06 PS=1.7e-06 $X=6855 $Y=2410 $dt=1
.ends HAJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DLY4JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DLY4JI3VX1 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=12 EP=4 FDC=12
M0 gnd3i! A 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.323e-13 AS=2.016e-13 PD=1.05e-06 PS=1.8e-06 $X=620 $Y=660 $dt=0
M1 8 10 gnd3i! gnd3i! ne3i L=1.8e-06 W=4.2e-07 AD=1.736e-13 AS=1.323e-13 PD=1.58e-06 PS=1.05e-06 $X=1600 $Y=660 $dt=0
M2 8 10 9 gnd3i! ne3i L=1.8e-06 W=4.2e-07 AD=1.736e-13 AS=2.00088e-13 PD=1.58e-06 PS=1.76778e-06 $X=1600 $Y=1360 $dt=0
M3 gnd3i! 9 7 gnd3i! ne3i L=1.1e-06 W=4.2e-07 AD=4.30324e-13 AS=2.16e-13 PD=1.75053e-06 PS=1.66e-06 $X=4630 $Y=660 $dt=0
M4 6 9 7 gnd3i! ne3i L=1.1e-06 W=4.2e-07 AD=2.00088e-13 AS=2.16e-13 PD=1.76778e-06 PS=1.66e-06 $X=4630 $Y=1400 $dt=0
M5 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.4055e-13 AS=9.11876e-13 PD=2.77e-06 PS=3.70947e-06 $X=7220 $Y=660 $dt=0
M6 vdd3i! A 10 vdd3i! pe3i L=3e-07 W=7e-07 AD=5.26875e-13 AS=3.535e-13 PD=3.30625e-06 PS=2.41e-06 $X=645 $Y=2680 $dt=1
M7 12 10 9 vdd3i! pe3i L=1.2e-06 W=4.2e-07 AD=1.674e-13 AS=2.016e-13 PD=1.56e-06 PS=1.8e-06 $X=2100 $Y=2680 $dt=1
M8 12 10 vdd3i! vdd3i! pe3i L=1.2e-06 W=4.2e-07 AD=1.674e-13 AS=3.16125e-13 PD=1.56e-06 PS=1.98375e-06 $X=2100 $Y=3400 $dt=1
M9 6 9 11 vdd3i! pe3i L=1.9e-06 W=4.2e-07 AD=2.016e-13 AS=1.674e-13 PD=1.8e-06 PS=1.56e-06 $X=4220 $Y=2680 $dt=1
M10 vdd3i! 9 11 vdd3i! pe3i L=1.9e-06 W=4.2e-07 AD=2.6367e-13 AS=1.674e-13 PD=1.32426e-06 PS=1.56e-06 $X=4220 $Y=3400 $dt=1
M11 Q 6 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.332e-13 AS=8.8518e-13 PD=3.86e-06 PS=4.44574e-06 $X=7245 $Y=2410 $dt=1
.ends DLY4JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO2I1JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO2I1JI3VX1 vdd3i! gnd3i! AN Q B
*.DEVICECLIMB
** N=8 EP=5 FDC=6
M0 gnd3i! AN 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.78131e-13 AS=2.016e-13 PD=1.19267e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 Q 7 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.4285e-13 AS=3.77469e-13 PD=1.445e-06 PS=2.52733e-06 $X=1460 $Y=660 $dt=0
M2 gnd3i! B Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=6.098e-13 AS=2.4285e-13 PD=3.52e-06 PS=1.445e-06 $X=2350 $Y=660 $dt=0
M3 vdd3i! AN 7 vdd3i! pe3i L=3e-07 W=7e-07 AD=4.32009e-13 AS=3.36e-13 PD=1.71185e-06 PS=2.36e-06 $X=620 $Y=2410 $dt=1
M4 8 7 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=8.70191e-13 PD=1.66e-06 PS=3.44815e-06 $X=1740 $Y=2410 $dt=1
M5 Q B 8 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=1.7625e-13 PD=3.78e-06 PS=1.66e-06 $X=2290 $Y=2410 $dt=1
.ends NO2I1JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AO22JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AO22JI3VX1 vdd3i! gnd3i! B A C D Q
*.DEVICECLIMB
** N=12 EP=7 FDC=10
M0 11 B gnd3i! gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=5.768e-13 PD=8.1e-07 PS=3.52e-06 $X=660 $Y=990 $dt=0
M1 10 A 11 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=1.68e-13 AS=7e-14 PD=1.16e-06 PS=8.1e-07 $X=1260 $Y=990 $dt=0
M2 9 C 10 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=1.68e-13 PD=8.1e-07 PS=1.16e-06 $X=2210 $Y=990 $dt=0
M3 gnd3i! D 9 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=3.96017e-13 AS=7e-14 PD=1.66069e-06 PS=8.1e-07 $X=2810 $Y=990 $dt=0
M4 Q 10 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=6.29383e-13 PD=2.74e-06 PS=2.63931e-06 $X=4070 $Y=660 $dt=0
M5 vdd3i! B 12 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=2.295e-13 AS=4.868e-13 PD=1.39e-06 PS=3.75e-06 $X=460 $Y=2490 $dt=1
M6 12 A vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.868e-13 AS=2.295e-13 PD=3.75e-06 PS=1.39e-06 $X=1300 $Y=2490 $dt=1
M7 10 C 12 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=2.295e-13 AS=4.868e-13 PD=1.39e-06 PS=3.75e-06 $X=2020 $Y=2490 $dt=1
M8 12 D 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.868e-13 AS=2.295e-13 PD=3.75e-06 PS=1.39e-06 $X=2860 $Y=2490 $dt=1
M9 Q 10 vdd3i! vdd3i! pe3i L=3.01705e-07 W=1.47627e-06 AD=5.312e-13 AS=7.778e-13 PD=3.68627e-06 PS=4.46627e-06 $X=4120 $Y=2410 $dt=1
.ends AO22JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX6                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX6 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=14
M0 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=6.008e-13 PD=1.34e-06 PS=3.52e-06 $X=660 $Y=750 $dt=0
M1 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=5.84805e-13 AS=2.16e-13 PD=2.17751e-06 PS=1.34e-06 $X=1550 $Y=750 $dt=0
M2 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=6.50595e-13 PD=1.43e-06 PS=2.42249e-06 $X=2960 $Y=660 $dt=0
M3 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=3850 $Y=660 $dt=0
M4 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=4820 $Y=660 $dt=0
M5 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=6.098e-13 AS=2.403e-13 PD=3.52e-06 PS=1.43e-06 $X=5710 $Y=660 $dt=0
M6 6 A vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=6.3285e-13 PD=1.87971e-06 PS=3.75971e-06 $X=525 $Y=2410 $dt=1
M7 vdd3i! A 6 vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=3.7905e-13 AS=2.751e-13 PD=1.98971e-06 PS=1.87971e-06 $X=1365 $Y=2410 $dt=1
M8 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=3.7905e-13 PD=1.87971e-06 PS=1.98971e-06 $X=2075 $Y=2410 $dt=1
M9 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=3.3675e-13 AS=2.751e-13 PD=1.92971e-06 PS=1.87971e-06 $X=2915 $Y=2410 $dt=1
M10 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=3.3675e-13 PD=1.87971e-06 PS=1.92971e-06 $X=3565 $Y=2410 $dt=1
M11 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=3.3675e-13 AS=2.751e-13 PD=1.92971e-06 PS=1.87971e-06 $X=4405 $Y=2410 $dt=1
M12 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=3.3675e-13 PD=1.87971e-06 PS=1.92971e-06 $X=5055 $Y=2410 $dt=1
M13 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=6.3285e-13 AS=2.751e-13 PD=3.75971e-06 PS=1.87971e-06 $X=5895 $Y=2410 $dt=1
.ends BUJI3VX6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ON31JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ON31JI3VX1 vdd3i! gnd3i! A B C Q D
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 9 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=6.098e-13 PD=1.43e-06 PS=3.52e-06 $X=660 $Y=660 $dt=0
M1 gnd3i! B 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=1550 $Y=660 $dt=0
M2 9 C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=2520 $Y=660 $dt=0
M3 Q D 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=2.403e-13 PD=2.74e-06 PS=1.43e-06 $X=3410 $Y=660 $dt=0
M4 11 A vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=9.066e-13 PD=1.72e-06 PS=4.59e-06 $X=1145 $Y=2410 $dt=1
M5 10 B 11 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=2.1855e-13 PD=1.72e-06 PS=1.72e-06 $X=1755 $Y=2410 $dt=1
M6 Q C 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=5.30442e-13 AS=2.1855e-13 PD=2.60067e-06 PS=1.72e-06 $X=2365 $Y=2410 $dt=1
M7 vdd3i! D Q vdd3i! pe3i L=3e-07 W=8.4e-07 AD=1.1576e-12 AS=3.16008e-13 PD=4.94e-06 PS=1.54933e-06 $X=3330 $Y=2410 $dt=1
.ends ON31JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: EO3JI3VX1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt EO3JI3VX1 vdd3i! gnd3i! C B A Q
*.DEVICECLIMB
** N=16 EP=6 FDC=20
M0 12 C gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.628e-13 PD=9.6e-07 PS=3.52e-06 $X=660 $Y=1130 $dt=0
M1 gnd3i! B 12 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.30196e-13 AS=1.134e-13 PD=1.36723e-06 PS=9.6e-07 $X=1550 $Y=1130 $dt=0
M2 11 C gnd3i! gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=6.5e-14 AS=2.85004e-13 PD=7.7e-07 PS=1.69277e-06 $X=2910 $Y=1030 $dt=0
M3 10 B 11 gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=1.404e-13 AS=6.5e-14 PD=1.06e-06 PS=7.7e-07 $X=3510 $Y=1030 $dt=0
M4 gnd3i! 12 10 gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=8.05779e-13 AS=1.404e-13 PD=2.83787e-06 PS=1.06e-06 $X=4400 $Y=1030 $dt=0
M5 9 10 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=6.50821e-13 PD=9.6e-07 PS=2.29213e-06 $X=6075 $Y=1130 $dt=0
M6 gnd3i! A 9 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.90537e-13 AS=1.134e-13 PD=1.53255e-06 PS=9.6e-07 $X=6965 $Y=1130 $dt=0
M7 8 A gnd3i! gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=6.5e-14 AS=3.59713e-13 PD=7.7e-07 PS=1.89745e-06 $X=8140 $Y=1030 $dt=0
M8 Q 10 8 gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=1.404e-13 AS=6.5e-14 PD=1.06e-06 PS=7.7e-07 $X=8740 $Y=1030 $dt=0
M9 gnd3i! 9 Q gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=5.728e-13 AS=1.404e-13 PD=3.52e-06 PS=1.06e-06 $X=9630 $Y=1030 $dt=0
M10 16 C vdd3i! vdd3i! pe3i L=3e-07 W=1.3e-06 AD=1.95e-13 AS=6.603e-13 PD=1.6e-06 PS=3.63e-06 $X=645 $Y=2520 $dt=1
M11 12 B 16 vdd3i! pe3i L=3e-07 W=1.3e-06 AD=5.157e-13 AS=1.95e-13 PD=3.61e-06 PS=1.6e-06 $X=1245 $Y=2520 $dt=1
M12 vdd3i! C 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=5.8645e-13 PD=2e-06 PS=3.83e-06 $X=2675 $Y=2410 $dt=1
M13 14 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=4.1595e-13 PD=2e-06 PS=2e-06 $X=3565 $Y=2410 $dt=1
M14 10 12 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=5.6965e-13 AS=4.1595e-13 PD=3.83e-06 PS=2e-06 $X=4455 $Y=2410 $dt=1
M15 15 10 vdd3i! vdd3i! pe3i L=3e-07 W=1.3e-06 AD=1.95e-13 AS=5.301e-13 PD=1.6e-06 PS=3.61e-06 $X=5885 $Y=2410 $dt=1
M16 9 A 15 vdd3i! pe3i L=3e-07 W=1.3e-06 AD=5.157e-13 AS=1.95e-13 PD=3.61e-06 PS=1.6e-06 $X=6485 $Y=2410 $dt=1
M17 vdd3i! A 13 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=5.8645e-13 PD=2e-06 PS=3.83e-06 $X=7915 $Y=2410 $dt=1
M18 13 10 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=4.1595e-13 PD=2e-06 PS=2e-06 $X=8805 $Y=2410 $dt=1
M19 Q 9 13 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.1205e-13 AS=4.1595e-13 PD=3.83e-06 PS=2e-06 $X=9695 $Y=2410 $dt=1
.ends EO3JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX2                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX2 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=6
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=6e-07 AD=2.96727e-13 AS=2.88e-13 PD=1.69091e-06 PS=2.16e-06 $X=620 $Y=950 $dt=0
M1 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=7.2e-07 AD=2.016e-13 AS=3.56073e-13 PD=1.512e-06 PS=2.02909e-06 $X=1590 $Y=830 $dt=0
M2 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=4.648e-13 AS=1.344e-13 PD=3.52e-06 PS=1.008e-06 $X=2480 $Y=1070 $dt=0
M3 vdd3i! A 6 vdd3i! pe3i L=3e-07 W=1.1e-06 AD=5.39943e-13 AS=5.28e-13 PD=2.20442e-06 PS=3.16e-06 $X=620 $Y=2410 $dt=1
M4 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=7.16507e-13 PD=1.87971e-06 PS=2.92528e-06 $X=1640 $Y=2410 $dt=1
M5 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=8.6265e-13 AS=2.751e-13 PD=4.56971e-06 PS=1.87971e-06 $X=2480 $Y=2410 $dt=1
.ends BUJI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INJI3VX3                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INJI3VX3 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=5 EP=4 FDC=5
M0 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=7.586e-13 PD=1.43e-06 PS=3.76e-06 $X=780 $Y=660 $dt=0
M1 gnd3i! A Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=7.586e-13 AS=2.403e-13 PD=3.76e-06 PS=1.43e-06 $X=1670 $Y=660 $dt=0
M2 Q A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=6.12287e-13 PD=1.86506e-06 PS=3.78506e-06 $X=490 $Y=2410 $dt=1
M3 vdd3i! A Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.86587e-13 AS=2.54913e-13 PD=1.88506e-06 PS=1.86506e-06 $X=1330 $Y=2410 $dt=1
M4 Q A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=5.51013e-13 AS=2.86587e-13 PD=3.69506e-06 PS=1.88506e-06 $X=1880 $Y=2410 $dt=1
.ends INJI3VX3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA3I2JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA3I2JI3VX1 vdd3i! gnd3i! AN BN C Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 9 AN gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=4.00432e-13 PD=9.6e-07 PS=2.10243e-06 $X=540 $Y=1130 $dt=0
M1 gnd3i! BN 9 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=4.00432e-13 AS=1.134e-13 PD=2.10243e-06 PS=9.6e-07 $X=1430 $Y=1130 $dt=0
M2 8 C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=8.48535e-13 PD=1.14e-06 PS=4.45514e-06 $X=2290 $Y=660 $dt=0
M3 Q 9 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.806e-13 AS=1.1125e-13 PD=2.86e-06 PS=1.14e-06 $X=2890 $Y=660 $dt=0
M4 10 AN 9 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=4.08e-13 PD=1.1e-06 PS=2.66e-06 $X=620 $Y=2410 $dt=1
M5 vdd3i! BN 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=7.38476e-13 AS=1.0625e-13 PD=3.31526e-06 PS=1.1e-06 $X=1170 $Y=2410 $dt=1
M6 vdd3i! C Q vdd3i! pe3i L=3.00037e-07 W=1.00071e-06 AD=8.69412e-13 AS=2.376e-13 PD=3.90308e-06 PS=1.49071e-06 $X=2170 $Y=2410 $dt=1
M7 Q 9 vdd3i! vdd3i! pe3i L=3.00037e-07 W=1.00071e-06 AD=2.376e-13 AS=8.69412e-13 PD=1.49071e-06 PS=3.90308e-06 $X=3010 $Y=2410 $dt=1
.ends NA3I2JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: EN3JI3VX1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt EN3JI3VX1 vdd3i! gnd3i! C B A Q
*.DEVICECLIMB
** N=16 EP=6 FDC=20
M0 13 C gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=2.016e-13 PD=9.6e-07 PS=1.8e-06 $X=620 $Y=1030 $dt=0
M1 gnd3i! B 13 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.97668e-13 AS=1.134e-13 PD=1.24213e-06 PS=9.6e-07 $X=1510 $Y=1030 $dt=0
M2 12 C gnd3i! gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=6.5e-14 AS=2.44732e-13 PD=7.7e-07 PS=1.53787e-06 $X=2730 $Y=930 $dt=0
M3 11 B 12 gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=1.404e-13 AS=6.5e-14 PD=1.06e-06 PS=7.7e-07 $X=3330 $Y=930 $dt=0
M4 gnd3i! 13 11 gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=5.308e-13 AS=1.404e-13 PD=3.32e-06 PS=1.06e-06 $X=4220 $Y=930 $dt=0
M5 9 11 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=5850 $Y=970 $dt=0
M6 gnd3i! A 9 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=6450 $Y=970 $dt=0
M7 8 A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=1.134e-13 PD=9.6e-07 PS=9.6e-07 $X=7340 $Y=970 $dt=0
M8 gnd3i! 11 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.965e-13 AS=1.134e-13 PD=3.17071e-06 PS=9.6e-07 $X=8230 $Y=970 $dt=0
M9 Q 10 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=2.0035e-13 PD=1.8e-06 PS=1.77071e-06 $X=9670 $Y=1130 $dt=0
M10 16 C vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.115e-13 AS=7.1585e-13 PD=1.71e-06 PS=3.85e-06 $X=645 $Y=2410 $dt=1
M11 13 B 16 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=5.5365e-13 AS=2.115e-13 PD=3.83e-06 PS=1.71e-06 $X=1245 $Y=2410 $dt=1
M12 vdd3i! C 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.23e-13 AS=5.8645e-13 PD=2.01e-06 PS=3.83e-06 $X=2675 $Y=2410 $dt=1
M13 14 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=4.23e-13 PD=2e-06 PS=2.01e-06 $X=3575 $Y=2410 $dt=1
M14 11 13 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.1205e-13 AS=4.1595e-13 PD=3.83e-06 PS=2e-06 $X=4465 $Y=2410 $dt=1
M15 10 11 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=9.1545e-13 PD=2e-06 PS=4.61e-06 $X=6095 $Y=2410 $dt=1
M16 vdd3i! A 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.956e-13 AS=4.1595e-13 PD=2.63e-06 PS=2e-06 $X=6985 $Y=2410 $dt=1
M17 15 A vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.115e-13 AS=6.956e-13 PD=1.71e-06 PS=2.63e-06 $X=8155 $Y=2410 $dt=1
M18 Q 11 15 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.66787e-13 AS=2.115e-13 PD=2.36668e-06 PS=1.71e-06 $X=8755 $Y=2410 $dt=1
M19 vdd3i! 10 Q vdd3i! pe3i L=3e-07 W=9.85e-07 AD=8.62325e-13 AS=3.26088e-13 PD=4.61e-06 PS=1.65332e-06 $X=9655 $Y=2410 $dt=1
.ends EN3JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: SDFRRQJI3VX1                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt SDFRRQJI3VX1 vdd3i! gnd3i! SE SD RN D C Q
*.DEVICECLIMB
** N=31 EP=8 FDC=39
M0 gnd3i! SE 25 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.11575e-13 AS=2.016e-13 PD=1.6275e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 13 RN gnd3i! gnd3i! ne3i L=3.5e-07 W=5.4e-07 AD=2.079e-13 AS=2.72025e-13 PD=1.4625e-06 PS=2.0925e-06 $X=1410 $Y=660 $dt=0
M2 24 SE 13 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.617e-13 PD=6.7e-07 PS=1.1375e-06 $X=2340 $Y=960 $dt=0
M3 12 SD 24 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.163e-13 AS=5.25e-14 PD=1.45e-06 PS=6.7e-07 $X=2940 $Y=960 $dt=0
M4 23 D 12 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.163e-13 PD=6.7e-07 PS=1.45e-06 $X=3910 $Y=1000 $dt=0
M5 13 25 23 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=5.25e-14 PD=1.8e-06 PS=6.7e-07 $X=4510 $Y=1000 $dt=0
M6 gnd3i! 20 22 gnd3i! ne3i L=3.5e-07 W=7.2e-07 AD=3.01862e-13 AS=3.456e-13 PD=1.65084e-06 PS=2.4e-06 $X=6100 $Y=1090 $dt=0
M7 11 RN gnd3i! gnd3i! ne3i L=3.5e-07 W=8.85e-07 AD=2.20538e-13 AS=3.71038e-13 PD=1.77e-06 PS=2.02916e-06 $X=7070 $Y=925 $dt=0
M8 21 22 11 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.04662e-13 PD=6.7e-07 PS=8.4e-07 $X=7840 $Y=1390 $dt=0
M9 20 18 21 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=8440 $Y=1390 $dt=0
M10 12 19 20 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=1.134e-13 PD=1.8e-06 PS=9.6e-07 $X=9330 $Y=1390 $dt=0
M11 gnd3i! C 19 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.722e-13 AS=2.016e-13 PD=1.24e-06 PS=1.8e-06 $X=10920 $Y=1390 $dt=0
M12 18 19 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=1.722e-13 PD=1.8e-06 PS=1.24e-06 $X=11930 $Y=1390 $dt=0
M13 17 22 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=13520 $Y=1020 $dt=0
M14 16 18 17 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=14120 $Y=1020 $dt=0
M15 15 19 16 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=15010 $Y=1020 $dt=0
M16 10 14 15 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.47785e-13 AS=5.25e-14 PD=9.42595e-07 PS=6.7e-07 $X=15610 $Y=1020 $dt=0
M17 gnd3i! RN 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.9815e-13 AS=3.13165e-13 PD=1.56e-06 PS=1.9974e-06 $X=16540 $Y=660 $dt=0
M18 14 16 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=2.9815e-13 PD=2.74e-06 PS=1.56e-06 $X=17560 $Y=660 $dt=0
M19 Q 16 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=6.098e-13 PD=2.74e-06 PS=3.52e-06 $X=19190 $Y=660 $dt=0
M20 vdd3i! SE 25 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=5.776e-13 AS=3.456e-13 PD=2.10667e-06 PS=2.4e-06 $X=620 $Y=2800 $dt=1
M21 31 25 vdd3i! vdd3i! pe3i L=3e-07 W=9e-07 AD=1.125e-13 AS=7.22e-13 PD=1.15e-06 PS=2.63333e-06 $X=2030 $Y=2620 $dt=1
M22 28 SD 31 vdd3i! pe3i L=3e-07 W=9e-07 AD=2.43e-13 AS=1.125e-13 PD=1.44e-06 PS=1.15e-06 $X=2580 $Y=2620 $dt=1
M23 30 D 28 vdd3i! pe3i L=3e-07 W=9e-07 AD=1.125e-13 AS=2.43e-13 PD=1.15e-06 PS=1.44e-06 $X=3420 $Y=2620 $dt=1
M24 vdd3i! SE 30 vdd3i! pe3i L=3e-07 W=9e-07 AD=3.80558e-13 AS=1.125e-13 PD=1.98274e-06 PS=1.15e-06 $X=3970 $Y=2620 $dt=1
M25 22 20 vdd3i! vdd3i! pe3i L=3e-07 W=1.07e-06 AD=5.136e-13 AS=4.52442e-13 PD=3.1e-06 PS=2.35726e-06 $X=4890 $Y=2745 $dt=1
M26 vdd3i! RN 20 vdd3i! pe3i L=3e-07 W=1.02e-06 AD=9.30148e-13 AS=4.896e-13 PD=3.58417e-06 PS=3e-06 $X=6430 $Y=2800 $dt=1
M27 29 22 vdd3i! vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=3.83002e-13 PD=6.7e-07 PS=1.47583e-06 $X=7890 $Y=3060 $dt=1
M28 20 19 29 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=1.218e-13 AS=5.25e-14 PD=9.22677e-07 PS=6.7e-07 $X=8440 $Y=3060 $dt=1
M29 28 18 20 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.08e-13 AS=2.465e-13 PD=2.66e-06 PS=1.86732e-06 $X=9285 $Y=2670 $dt=1
M30 19 C vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.0675e-13 AS=6.327e-13 PD=2.37071e-06 PS=3.56e-06 $X=10970 $Y=2735 $dt=1
M31 vdd3i! 19 18 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.27981e-13 AS=4.01587e-13 PD=1.59258e-06 PS=3.03778e-06 $X=12390 $Y=2800 $dt=1
M32 27 22 vdd3i! vdd3i! pe3i L=3e-07 W=7.9e-07 AD=1.16525e-13 AS=3.59869e-13 PD=1.085e-06 PS=1.74742e-06 $X=13570 $Y=2730 $dt=1
M33 16 19 27 vdd3i! pe3i L=3e-07 W=7.9e-07 AD=2.25379e-13 AS=1.16525e-13 PD=1.73669e-06 PS=1.085e-06 $X=14165 $Y=2730 $dt=1
M34 26 18 16 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=1.19821e-13 PD=6.7e-07 PS=9.23306e-07 $X=15005 $Y=3100 $dt=1
M35 vdd3i! 14 26 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=6.29844e-13 AS=5.25e-14 PD=2.86017e-06 PS=6.7e-07 $X=15555 $Y=3100 $dt=1
M36 vdd3i! RN 16 vdd3i! pe3i L=3e-07 W=7.9e-07 AD=1.18471e-12 AS=3.19387e-13 PD=5.37983e-06 PS=2.5195e-06 $X=16775 $Y=2410 $dt=1
M37 vdd3i! 16 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=6.768e-13 PD=1.95e-06 PS=3.78e-06 $X=18400 $Y=2410 $dt=1
M38 Q 16 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=3.807e-13 PD=3.78e-06 PS=1.95e-06 $X=19240 $Y=2410 $dt=1
.ends SDFRRQJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO2JI3VX0 vdd3i! gnd3i! B Q A
*.DEVICECLIMB
** N=7 EP=5 FDC=4
M0 Q B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=7.244e-13 PD=9.6e-07 PS=4.14e-06 $X=500 $Y=1130 $dt=0
M1 gnd3i! A Q gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=7.244e-13 AS=1.134e-13 PD=4.14e-06 PS=9.6e-07 $X=1390 $Y=1130 $dt=0
M2 7 B vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=9.298e-13 PD=1.1e-06 PS=4.68e-06 $X=720 $Y=2410 $dt=1
M3 Q A 7 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.08e-13 AS=1.0625e-13 PD=2.66e-06 PS=1.1e-06 $X=1270 $Y=2410 $dt=1
.ends NO2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA4JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA4JI3VX0 vdd3i! gnd3i! D Q C B A
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 11 D gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=1.2e-13 AS=7.868e-13 PD=1.1e-06 PS=3.82e-06 $X=810 $Y=750 $dt=0
M1 10 C 11 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=1.2e-13 AS=1.2e-13 PD=1.1e-06 PS=1.1e-06 $X=1460 $Y=750 $dt=0
M2 9 B 10 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=1.2e-13 AS=1.2e-13 PD=1.1e-06 PS=1.1e-06 $X=2110 $Y=750 $dt=0
M3 Q A 9 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.84e-13 AS=1.2e-13 PD=2.56e-06 PS=1.1e-06 $X=2760 $Y=750 $dt=0
M4 Q D vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=9.882e-13 PD=1.24e-06 PS=3.92e-06 $X=540 $Y=2410 $dt=1
M5 vdd3i! C Q vdd3i! pe3i L=3e-07 W=7e-07 AD=9.882e-13 AS=1.89e-13 PD=3.92e-06 PS=1.24e-06 $X=1380 $Y=2410 $dt=1
M6 Q B vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=9.882e-13 PD=1.24e-06 PS=3.92e-06 $X=2240 $Y=2410 $dt=1
M7 vdd3i! A Q vdd3i! pe3i L=3e-07 W=7e-07 AD=9.882e-13 AS=1.89e-13 PD=3.92e-06 PS=1.24e-06 $X=3080 $Y=2410 $dt=1
.ends NA4JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA2JI3VX0 vdd3i! gnd3i! B Q A
*.DEVICECLIMB
** N=7 EP=5 FDC=4
M0 7 B gnd3i! gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=5.892e-13 PD=8.1e-07 PS=3.54e-06 $X=670 $Y=990 $dt=0
M1 Q A 7 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=2.688e-13 AS=7e-14 PD=2.08e-06 PS=8.1e-07 $X=1270 $Y=990 $dt=0
M2 Q B vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=1.1114e-12 PD=1.24e-06 PS=4.94e-06 $X=550 $Y=2410 $dt=1
M3 vdd3i! A Q vdd3i! pe3i L=3e-07 W=7e-07 AD=1.1114e-12 AS=1.89e-13 PD=4.94e-06 PS=1.24e-06 $X=1390 $Y=2410 $dt=1
.ends NA2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ON21JI3VX4                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ON21JI3VX4 vdd3i! gnd3i! B A C Q
*.DEVICECLIMB
** N=11 EP=6 FDC=16
M0 gnd3i! B 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=4.272e-13 PD=1.43e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 10 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=1510 $Y=660 $dt=0
M2 9 C 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.868e-13 AS=2.403e-13 PD=2.70971e-06 PS=1.43e-06 $X=2400 $Y=660 $dt=0
M3 gnd3i! 9 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.35783e-13 AS=4.34e-13 PD=1.42065e-06 PS=2.92971e-06 $X=3930 $Y=660 $dt=0
M4 Q 8 gnd3i! gnd3i! ne3i L=3.49164e-07 W=8.96213e-07 AD=2.32912e-13 AS=2.37429e-13 PD=1.42121e-06 PS=1.43057e-06 $X=4820 $Y=660 $dt=0
M5 gnd3i! 8 Q gnd3i! ne3i L=3.49164e-07 W=8.96213e-07 AD=2.32912e-13 AS=2.32912e-13 PD=1.42121e-06 PS=1.42121e-06 $X=5680 $Y=660 $dt=0
M6 Q 8 gnd3i! gnd3i! ne3i L=3.49164e-07 W=8.96213e-07 AD=2.32912e-13 AS=2.32912e-13 PD=1.42121e-06 PS=1.42121e-06 $X=6570 $Y=660 $dt=0
M7 gnd3i! 8 Q gnd3i! ne3i L=3.49164e-07 W=8.96213e-07 AD=4.19812e-13 AS=2.32912e-13 PD=2.73121e-06 PS=1.42121e-06 $X=7430 $Y=660 $dt=0
M8 11 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=9.418e-13 PD=1.66e-06 PS=4.63e-06 $X=695 $Y=2410 $dt=1
M9 9 A 11 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.68825e-13 AS=1.7625e-13 PD=2.075e-06 PS=1.66e-06 $X=1245 $Y=2410 $dt=1
M10 vdd3i! C 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.285e-12 AS=4.68825e-13 PD=5.02e-06 PS=2.075e-06 $X=2210 $Y=2410 $dt=1
M11 vdd3i! 9 8 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=5.48179e-13 AS=6.768e-13 PD=2.4141e-06 PS=3.78e-06 $X=4020 $Y=2410 $dt=1
M12 Q 8 vdd3i! vdd3i! pe3i L=3.00021e-07 W=1.42657e-06 AD=3.433e-13 AS=5.54621e-13 PD=1.92657e-06 PS=2.44247e-06 $X=4960 $Y=2410 $dt=1
M13 vdd3i! 8 Q vdd3i! pe3i L=3.00021e-07 W=1.42657e-06 AD=4.866e-13 AS=3.433e-13 PD=2.35657e-06 PS=1.92657e-06 $X=5800 $Y=2410 $dt=1
M14 Q 8 vdd3i! vdd3i! pe3i L=3.00021e-07 W=1.42657e-06 AD=3.433e-13 AS=4.866e-13 PD=1.92657e-06 PS=2.35657e-06 $X=6640 $Y=2410 $dt=1
M15 vdd3i! 8 Q vdd3i! pe3i L=3.00021e-07 W=1.42657e-06 AD=8.562e-13 AS=3.433e-13 PD=4.53657e-06 PS=1.92657e-06 $X=7480 $Y=2410 $dt=1
.ends ON21JI3VX4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND2JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND2JI3VX1 vdd3i! gnd3i! A B Q
*.DEVICECLIMB
** N=8 EP=5 FDC=6
M0 7 A 8 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=2.688e-13 PD=8.1e-07 PS=2.08e-06 $X=820 $Y=990 $dt=0
M1 gnd3i! B 7 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=2.57137e-13 AS=7e-14 PD=1.43669e-06 PS=8.1e-07 $X=1420 $Y=990 $dt=0
M2 Q 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=4.08663e-13 PD=2.74e-06 PS=2.28331e-06 $X=2390 $Y=660 $dt=0
M3 8 A vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=7.276e-13 PD=1.24e-06 PS=4.56e-06 $X=580 $Y=2410 $dt=1
M4 vdd3i! B 8 vdd3i! pe3i L=3e-07 W=7e-07 AD=3.64829e-13 AS=1.89e-13 PD=1.6455e-06 PS=1.24e-06 $X=1420 $Y=2410 $dt=1
M5 Q 8 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=7.34871e-13 PD=3.78e-06 PS=3.3145e-06 $X=2440 $Y=2410 $dt=1
.ends AND2JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA4JI3VX2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA4JI3VX2 vdd3i! gnd3i! Q D C B A
*.DEVICECLIMB
** N=14 EP=7 FDC=16
M0 14 D gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.78e-13 AS=6.098e-13 PD=1.29e-06 PS=3.52e-06 $X=660 $Y=660 $dt=0
M1 13 C 14 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.8245e-13 AS=1.78e-13 PD=1.3e-06 PS=1.29e-06 $X=1410 $Y=660 $dt=0
M2 12 B 13 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.78e-13 AS=1.8245e-13 PD=1.29e-06 PS=1.3e-06 $X=2170 $Y=660 $dt=0
M3 Q A 12 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.293e-13 AS=1.78e-13 PD=1.63e-06 PS=1.29e-06 $X=2920 $Y=660 $dt=0
M4 11 A Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.78e-13 AS=3.293e-13 PD=1.29e-06 PS=1.63e-06 $X=4010 $Y=660 $dt=0
M5 10 B 11 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.8245e-13 AS=1.78e-13 PD=1.3e-06 PS=1.29e-06 $X=4760 $Y=660 $dt=0
M6 9 C 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.78e-13 AS=1.8245e-13 PD=1.29e-06 PS=1.3e-06 $X=5520 $Y=660 $dt=0
M7 gnd3i! D 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=6.098e-13 AS=1.78e-13 PD=3.52e-06 PS=1.29e-06 $X=6270 $Y=660 $dt=0
M8 vdd3i! D Q vdd3i! pe3i L=3.00056e-07 W=9.91066e-07 AD=6.12287e-13 AS=4.22737e-13 PD=2.90357e-06 PS=2.83607e-06 $X=620 $Y=2410 $dt=1
M9 vdd3i! C Q vdd3i! pe3i L=3.00056e-07 W=9.91066e-07 AD=6.12287e-13 AS=2.21137e-13 PD=2.90357e-06 PS=1.45607e-06 $X=1440 $Y=2410 $dt=1
M10 Q B vdd3i! vdd3i! pe3i L=3.00056e-07 W=9.91066e-07 AD=2.21137e-13 AS=6.12287e-13 PD=1.45607e-06 PS=2.90357e-06 $X=2280 $Y=2410 $dt=1
M11 vdd3i! A Q vdd3i! pe3i L=3.00056e-07 W=9.91066e-07 AD=6.12287e-13 AS=2.93137e-13 PD=2.90357e-06 PS=1.60607e-06 $X=2995 $Y=2410 $dt=1
M12 Q A vdd3i! vdd3i! pe3i L=3.00056e-07 W=9.91066e-07 AD=2.93137e-13 AS=6.12287e-13 PD=1.60607e-06 PS=2.90357e-06 $X=3985 $Y=2410 $dt=1
M13 vdd3i! B Q vdd3i! pe3i L=3.00056e-07 W=9.91066e-07 AD=6.12287e-13 AS=2.21137e-13 PD=2.90357e-06 PS=1.45607e-06 $X=4700 $Y=2410 $dt=1
M14 Q C vdd3i! vdd3i! pe3i L=3.00056e-07 W=9.91066e-07 AD=2.21137e-13 AS=6.12287e-13 PD=1.45607e-06 PS=2.90357e-06 $X=5540 $Y=2410 $dt=1
M15 Q D vdd3i! vdd3i! pe3i L=3.00056e-07 W=9.91066e-07 AD=4.22737e-13 AS=6.12287e-13 PD=2.83607e-06 PS=2.90357e-06 $X=6360 $Y=2410 $dt=1
.ends NA4JI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO2I1JI3VX2                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO2I1JI3VX2 vdd3i! gnd3i! AN Q B
*.DEVICECLIMB
** N=9 EP=5 FDC=10
M0 gnd3i! AN 7 gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.3695e-13 AS=4.15012e-13 PD=1.44536e-06 PS=2.72536e-06 $X=595 $Y=660 $dt=0
M1 Q 7 gnd3i! gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.28113e-13 AS=2.3695e-13 PD=1.41536e-06 PS=1.44536e-06 $X=1500 $Y=660 $dt=0
M2 gnd3i! B Q gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.30162e-13 AS=2.28113e-13 PD=1.43036e-06 PS=1.41536e-06 $X=2340 $Y=660 $dt=0
M3 Q B gnd3i! gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.28113e-13 AS=2.30162e-13 PD=1.41536e-06 PS=1.43036e-06 $X=3230 $Y=660 $dt=0
M4 gnd3i! 7 Q gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=4.20212e-13 AS=2.28113e-13 PD=2.75536e-06 PS=1.41536e-06 $X=4070 $Y=660 $dt=0
M5 vdd3i! AN 7 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.998e-13 AS=6.768e-13 PD=2.595e-06 PS=3.78e-06 $X=620 $Y=2410 $dt=1
M6 9 7 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.115e-13 AS=6.998e-13 PD=1.71e-06 PS=2.595e-06 $X=1755 $Y=2410 $dt=1
M7 Q B 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.8775e-13 AS=2.115e-13 PD=1.96e-06 PS=1.71e-06 $X=2355 $Y=2410 $dt=1
M8 8 B Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.115e-13 AS=3.8775e-13 PD=1.71e-06 PS=1.96e-06 $X=3205 $Y=2410 $dt=1
M9 vdd3i! 7 8 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.3642e-12 AS=2.115e-13 PD=5.11e-06 PS=1.71e-06 $X=3805 $Y=2410 $dt=1
.ends NO2I1JI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: EO2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt EO2JI3VX0 vdd3i! gnd3i! B A Q
*.DEVICECLIMB
** N=10 EP=5 FDC=10
M0 8 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.628e-13 PD=9.6e-07 PS=3.52e-06 $X=660 $Y=1130 $dt=0
M1 gnd3i! A 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.0445e-13 AS=1.134e-13 PD=1.34e-06 PS=9.6e-07 $X=1550 $Y=1130 $dt=0
M2 7 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.0445e-13 PD=6.7e-07 PS=1.34e-06 $X=2670 $Y=980 $dt=0
M3 Q A 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.503e-13 AS=5.25e-14 PD=1.15e-06 PS=6.7e-07 $X=3270 $Y=980 $dt=0
M4 gnd3i! 8 Q gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.0464e-12 AS=1.503e-13 PD=4.3e-06 PS=1.15e-06 $X=4200 $Y=1130 $dt=0
M5 10 B vdd3i! vdd3i! pe3i L=3e-07 W=9e-07 AD=1.35e-13 AS=7.175e-13 PD=1.2e-06 PS=4.61e-06 $X=575 $Y=2410 $dt=1
M6 8 A 10 vdd3i! pe3i L=3e-07 W=9e-07 AD=5.38188e-13 AS=1.35e-13 PD=3.13778e-06 PS=1.2e-06 $X=1175 $Y=2410 $dt=1
M7 vdd3i! B 9 vdd3i! pe3i L=3e-07 W=1.3e-06 AD=5.321e-13 AS=5.76588e-13 PD=2.43e-06 PS=3.57778e-06 $X=2795 $Y=2520 $dt=1
M8 9 A vdd3i! vdd3i! pe3i L=3e-07 W=1.3e-06 AD=3.835e-13 AS=5.321e-13 PD=1.89e-06 PS=2.43e-06 $X=3765 $Y=2410 $dt=1
M9 Q 8 9 vdd3i! pe3i L=3e-07 W=1.3e-06 AD=6.565e-13 AS=3.835e-13 PD=3.61e-06 PS=1.89e-06 $X=4655 $Y=2410 $dt=1
.ends EO2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND2JI3VX0                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND2JI3VX0 vdd3i! gnd3i! A B Q
*.DEVICECLIMB
** N=8 EP=5 FDC=6
M0 7 A 8 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=2.688e-13 PD=8.1e-07 PS=2.08e-06 $X=820 $Y=990 $dt=0
M1 gnd3i! B 7 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=3.536e-13 AS=7e-14 PD=2.12571e-06 PS=8.1e-07 $X=1420 $Y=990 $dt=0
M2 Q 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=2.652e-13 PD=1.8e-06 PS=1.59429e-06 $X=2390 $Y=1130 $dt=0
M3 8 A vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=7.276e-13 PD=1.24e-06 PS=4.56e-06 $X=580 $Y=2410 $dt=1
M4 vdd3i! B 8 vdd3i! pe3i L=3e-07 W=7e-07 AD=5.276e-13 AS=1.89e-13 PD=2.48e-06 PS=1.24e-06 $X=1420 $Y=2410 $dt=1
M5 Q 8 vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=3.36e-13 AS=5.276e-13 PD=2.36e-06 PS=2.48e-06 $X=2440 $Y=2410 $dt=1
.ends AND2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AN22JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AN22JI3VX1 vdd3i! gnd3i! B A Q C D
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 10 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=6.098e-13 PD=1.14e-06 PS=3.52e-06 $X=660 $Y=660 $dt=0
M1 Q A 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=1.1125e-13 PD=1.43e-06 PS=1.14e-06 $X=1260 $Y=660 $dt=0
M2 9 C Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=2.403e-13 PD=1.14e-06 PS=1.43e-06 $X=2150 $Y=660 $dt=0
M3 gnd3i! D 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=8.082e-13 AS=1.1125e-13 PD=3.84e-06 PS=1.14e-06 $X=2750 $Y=660 $dt=0
M4 vdd3i! B 11 vdd3i! pe3i L=3.01094e-07 W=1.47213e-06 AD=4.29e-13 AS=6.0945e-13 PD=2.32213e-06 PS=3.77213e-06 $X=660 $Y=2410 $dt=1
M5 11 A vdd3i! vdd3i! pe3i L=3.01094e-07 W=1.47213e-06 AD=4.05825e-13 AS=4.29e-13 PD=2.06213e-06 PS=2.32213e-06 $X=1310 $Y=2410 $dt=1
M6 Q C 11 vdd3i! pe3i L=3.01094e-07 W=1.47213e-06 AD=2.9925e-13 AS=4.05825e-13 PD=1.92213e-06 PS=2.06213e-06 $X=2200 $Y=2410 $dt=1
M7 11 D Q vdd3i! pe3i L=3.01094e-07 W=1.47213e-06 AD=6.252e-13 AS=2.9925e-13 PD=3.77213e-06 PS=1.92213e-06 $X=3100 $Y=2410 $dt=1
.ends AN22JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO2JI3VX2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO2JI3VX2 vdd3i! gnd3i! B A Q
*.DEVICECLIMB
** N=8 EP=5 FDC=8
M0 Q B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=6.842e-13 PD=1.43e-06 PS=3.64e-06 $X=720 $Y=660 $dt=0
M1 gnd3i! A Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=1610 $Y=660 $dt=0
M2 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=2580 $Y=660 $dt=0
M3 gnd3i! B Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=6.098e-13 AS=2.403e-13 PD=3.52e-06 PS=1.43e-06 $X=3470 $Y=660 $dt=0
M4 8 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=1.6898e-12 PD=1.66e-06 PS=5.48e-06 $X=1120 $Y=2410 $dt=1
M5 Q A 8 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=1.7625e-13 PD=1.95e-06 PS=1.66e-06 $X=1670 $Y=2410 $dt=1
M6 7 A Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=3.807e-13 PD=1.66e-06 PS=1.95e-06 $X=2510 $Y=2410 $dt=1
M7 vdd3i! B 7 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.6898e-12 AS=1.7625e-13 PD=5.48e-06 PS=1.66e-06 $X=3060 $Y=2410 $dt=1
.ends NO2JI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AO21JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AO21JI3VX1 vdd3i! gnd3i! B A C Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 9 B gnd3i! gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=5.768e-13 PD=8.1e-07 PS=3.52e-06 $X=660 $Y=990 $dt=0
M1 8 A 9 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=1.708e-13 AS=7e-14 PD=1.17e-06 PS=8.1e-07 $X=1260 $Y=990 $dt=0
M2 gnd3i! C 8 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=3.94626e-13 AS=1.708e-13 PD=1.68386e-06 PS=1.17e-06 $X=2220 $Y=990 $dt=0
M3 Q 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=6.27174e-13 PD=2.74e-06 PS=2.67614e-06 $X=3510 $Y=660 $dt=0
M4 vdd3i! B 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=3.8185e-13 AS=4.08e-13 PD=2.53e-06 PS=2.66e-06 $X=620 $Y=2410 $dt=1
M5 10 A vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=2.295e-13 AS=3.8185e-13 PD=1.39e-06 PS=2.53e-06 $X=1340 $Y=2410 $dt=1
M6 8 C 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.08e-13 AS=2.295e-13 PD=2.66e-06 PS=1.39e-06 $X=2180 $Y=2410 $dt=1
M7 Q 8 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=7.0775e-13 PD=3.78e-06 PS=4.73e-06 $X=3560 $Y=2410 $dt=1
.ends AO21JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA2I1JI3VX2                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA2I1JI3VX2 vdd3i! gnd3i! AN Q B
*.DEVICECLIMB
** N=9 EP=5 FDC=10
M0 gnd3i! AN 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.672e-13 AS=4.272e-13 PD=2.05e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 8 9 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=4.672e-13 PD=1.14e-06 PS=2.05e-06 $X=1780 $Y=660 $dt=0
M2 Q B 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.759e-13 AS=1.1125e-13 PD=1.51e-06 PS=1.14e-06 $X=2380 $Y=660 $dt=0
M3 7 B Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=2.759e-13 PD=1.14e-06 PS=1.51e-06 $X=3350 $Y=660 $dt=0
M4 gnd3i! 9 7 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=7.09e-13 AS=1.1125e-13 PD=3.68e-06 PS=1.14e-06 $X=3950 $Y=660 $dt=0
M5 vdd3i! AN 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=9.9878e-13 AS=6.768e-13 PD=4.57664e-06 PS=3.78e-06 $X=620 $Y=2410 $dt=1
M6 Q 9 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.7e-13 AS=7.08355e-13 PD=1.54e-06 PS=3.24584e-06 $X=1540 $Y=2410 $dt=1
M7 vdd3i! B Q vdd3i! pe3i L=3e-07 W=1e-06 AD=7.08355e-13 AS=2.7e-13 PD=3.24584e-06 PS=1.54e-06 $X=2380 $Y=2410 $dt=1
M8 Q B vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.7e-13 AS=7.08355e-13 PD=1.54e-06 PS=3.24584e-06 $X=3280 $Y=2410 $dt=1
M9 vdd3i! 9 Q vdd3i! pe3i L=3e-07 W=1e-06 AD=7.08355e-13 AS=2.7e-13 PD=3.24584e-06 PS=1.54e-06 $X=4120 $Y=2410 $dt=1
.ends NA2I1JI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA22JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA22JI3VX1 vdd3i! gnd3i! A B C Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 9 A 10 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=2.688e-13 PD=8.1e-07 PS=2.08e-06 $X=620 $Y=990 $dt=0
M1 gnd3i! B 9 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=3.3376e-13 AS=7e-14 PD=1.56028e-06 PS=8.1e-07 $X=1220 $Y=990 $dt=0
M2 8 C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=5.3044e-13 PD=1.14e-06 PS=2.47972e-06 $X=2350 $Y=660 $dt=0
M3 Q 10 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=1.1125e-13 PD=2.74e-06 PS=1.14e-06 $X=2950 $Y=660 $dt=0
M4 10 A vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=7.66562e-13 PD=1.24e-06 PS=3.33273e-06 $X=510 $Y=2410 $dt=1
M5 vdd3i! B 10 vdd3i! pe3i L=3e-07 W=7e-07 AD=7.66562e-13 AS=1.89e-13 PD=3.33273e-06 PS=1.24e-06 $X=1350 $Y=2410 $dt=1
M6 vdd3i! C Q vdd3i! pe3i L=3.00052e-07 W=9.98995e-07 AD=1.09399e-12 AS=2.255e-13 PD=4.75626e-06 PS=1.46899e-06 $X=2190 $Y=2410 $dt=1
M7 Q 10 vdd3i! vdd3i! pe3i L=3.00052e-07 W=9.98995e-07 AD=2.255e-13 AS=1.09399e-12 PD=1.46899e-06 PS=4.75626e-06 $X=3030 $Y=2410 $dt=1
.ends NA22JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MU2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MU2JI3VX0 vdd3i! gnd3i! S IN0 IN1 Q
*.DEVICECLIMB
** N=13 EP=6 FDC=12
M0 gnd3i! S 11 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.5315e-13 AS=2.016e-13 PD=1.165e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 10 IN0 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.5315e-13 PD=6.7e-07 PS=1.165e-06 $X=1550 $Y=965 $dt=0
M2 9 11 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=2150 $Y=965 $dt=0
M3 8 S 9 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=3040 $Y=965 $dt=0
M4 gnd3i! IN1 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.148e-13 AS=5.25e-14 PD=1.88e-06 PS=6.7e-07 $X=3640 $Y=965 $dt=0
M5 Q 9 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=3.148e-13 PD=1.8e-06 PS=1.88e-06 $X=4630 $Y=1130 $dt=0
M6 vdd3i! S 11 vdd3i! pe3i L=3e-07 W=5e-07 AD=1.78281e-13 AS=2.525e-13 PD=1.10156e-06 PS=2.01e-06 $X=645 $Y=2675 $dt=1
M7 13 IN0 vdd3i! vdd3i! pe3i L=3e-07 W=7.8e-07 AD=1.17e-13 AS=2.78119e-13 PD=1.08e-06 PS=1.71844e-06 $X=1575 $Y=2675 $dt=1
M8 9 S 13 vdd3i! pe3i L=3e-07 W=7.8e-07 AD=2.301e-13 AS=1.17e-13 PD=1.37e-06 PS=1.08e-06 $X=2175 $Y=2675 $dt=1
M9 12 11 9 vdd3i! pe3i L=3e-07 W=7.8e-07 AD=1.17e-13 AS=2.301e-13 PD=1.08e-06 PS=1.37e-06 $X=3065 $Y=2675 $dt=1
M10 vdd3i! IN1 12 vdd3i! pe3i L=3e-07 W=7.8e-07 AD=5.0563e-13 AS=1.17e-13 PD=2.58243e-06 PS=1.08e-06 $X=3665 $Y=2675 $dt=1
M11 Q 9 vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=3.535e-13 AS=4.5377e-13 PD=2.41e-06 PS=2.31757e-06 $X=4655 $Y=2410 $dt=1
.ends MU2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OR3JI3VX1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OR3JI3VX1 vdd3i! gnd3i! A B C Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 gnd3i! A 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.482e-13 AS=2.016e-13 PD=2.04e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 8 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.116e-13 AS=2.482e-13 PD=1.78e-06 PS=2.04e-06 $X=1390 $Y=1310 $dt=0
M2 gnd3i! C 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.66689e-13 AS=2.116e-13 PD=1.17398e-06 PS=1.78e-06 $X=2160 $Y=1130 $dt=0
M3 Q 8 gnd3i! gnd3i! ne3i L=3.50112e-07 W=8.98284e-07 AD=4.174e-13 AS=3.56511e-13 PD=2.72828e-06 PS=2.51087e-06 $X=2970 $Y=660 $dt=0
M4 10 A 8 vdd3i! pe3i L=3e-07 W=1e-06 AD=1.375e-13 AS=4.8e-13 PD=1.275e-06 PS=2.96e-06 $X=670 $Y=2720 $dt=1
M5 9 B 10 vdd3i! pe3i L=3e-07 W=1e-06 AD=1.375e-13 AS=1.375e-13 PD=1.275e-06 PS=1.275e-06 $X=1245 $Y=2720 $dt=1
M6 vdd3i! C 9 vdd3i! pe3i L=3e-07 W=1e-06 AD=5.59502e-13 AS=1.375e-13 PD=2.19087e-06 PS=1.275e-06 $X=1820 $Y=2720 $dt=1
M7 Q 8 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=7.88898e-13 PD=3.78e-06 PS=3.08913e-06 $X=3000 $Y=2410 $dt=1
.ends OR3JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ON211JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ON211JI3VX1 vdd3i! gnd3i! B Q A C D
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 Q B 10 gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.27987e-13 AS=4.20337e-13 PD=1.41536e-06 PS=2.75536e-06 $X=620 $Y=660 $dt=0
M1 10 A Q gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.30287e-13 AS=2.27987e-13 PD=1.43036e-06 PS=1.41536e-06 $X=1460 $Y=660 $dt=0
M2 9 C 10 gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=1.21188e-13 AS=2.30287e-13 PD=1.17536e-06 PS=1.43036e-06 $X=2350 $Y=660 $dt=0
M3 gnd3i! D 9 gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=4.20337e-13 AS=1.21188e-13 PD=2.75536e-06 PS=1.17536e-06 $X=2950 $Y=660 $dt=0
M4 11 B vdd3i! vdd3i! pe3i L=3e-07 W=1.38e-06 AD=1.725e-13 AS=9.388e-13 PD=1.63e-06 PS=4.63e-06 $X=695 $Y=2410 $dt=1
M5 Q A 11 vdd3i! pe3i L=3e-07 W=1.38e-06 AD=4.69617e-13 AS=1.725e-13 PD=2.38255e-06 PS=1.63e-06 $X=1245 $Y=2410 $dt=1
M6 vdd3i! C Q vdd3i! pe3i L=3.00049e-07 W=9.66924e-07 AD=4.25413e-13 AS=3.29046e-13 PD=2.34192e-06 PS=1.66938e-06 $X=2210 $Y=2410 $dt=1
M7 Q D vdd3i! vdd3i! pe3i L=3.00049e-07 W=9.66924e-07 AD=4.20162e-13 AS=4.25413e-13 PD=2.80192e-06 PS=2.34192e-06 $X=3000 $Y=2410 $dt=1
.ends ON211JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AN21JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AN21JI3VX1 vdd3i! gnd3i! B A Q C
*.DEVICECLIMB
** N=9 EP=6 FDC=6
M0 8 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=6.47e-13 PD=1.14e-06 PS=3.58e-06 $X=690 $Y=660 $dt=0
M1 Q A 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.28413e-13 AS=1.1125e-13 PD=1.78572e-06 PS=1.14e-06 $X=1290 $Y=660 $dt=0
M2 gnd3i! C Q gnd3i! ne3i L=3.5e-07 W=6.65e-07 AD=6.369e-13 AS=2.45387e-13 PD=3.6e-06 PS=1.33428e-06 $X=2310 $Y=885 $dt=0
M3 vdd3i! B 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.371e-13 AS=6.768e-13 PD=2.03e-06 PS=3.78e-06 $X=620 $Y=2410 $dt=1
M4 9 A vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=4.371e-13 PD=1.95e-06 PS=2.03e-06 $X=1540 $Y=2410 $dt=1
M5 Q C 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.614e-13 AS=3.807e-13 PD=3.9e-06 PS=1.95e-06 $X=2380 $Y=2410 $dt=1
.ends AN21JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INJI3VX0                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INJI3VX0 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=5 EP=4 FDC=2
M0 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=6.248e-13 PD=1.8e-06 PS=3.62e-06 $X=710 $Y=1130 $dt=0
M1 Q A vdd3i! vdd3i! pe3i L=3e-07 W=9.4e-07 AD=4.512e-13 AS=1.0092e-12 PD=2.84e-06 PS=4.76e-06 $X=760 $Y=2410 $dt=1
.ends INJI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO3I1JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO3I1JI3VX1 vdd3i! gnd3i! AN Q B C
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 gnd3i! AN 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.99484e-13 AS=2.016e-13 PD=1.19267e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 Q 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=4.22716e-13 PD=1.43e-06 PS=2.52733e-06 $X=1550 $Y=660 $dt=0
M2 gnd3i! B Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=2440 $Y=660 $dt=0
M3 Q C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=3.494e-13 PD=2.74e-06 PS=1.86e-06 $X=3410 $Y=660 $dt=0
M4 vdd3i! AN 8 vdd3i! pe3i L=3e-07 W=7e-07 AD=4.49443e-13 AS=3.36e-13 PD=1.73175e-06 PS=2.36e-06 $X=620 $Y=2415 $dt=1
M5 10 8 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=9.05307e-13 PD=1.72e-06 PS=3.48825e-06 $X=1770 $Y=2410 $dt=1
M6 9 B 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=2.1855e-13 PD=1.72e-06 PS=1.72e-06 $X=2380 $Y=2410 $dt=1
M7 Q C 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=2.1855e-13 PD=3.78e-06 PS=1.72e-06 $X=2990 $Y=2410 $dt=1
.ends NO3I1JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP25JI3V                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP25JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=12
M0 gnd3i! 5 4 gnd3i! ne3i L=3.5e-07 W=8.8e-07 AD=2.376e-13 AS=4.224e-13 PD=1.42e-06 PS=2.72e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=1510 $Y=660 $dt=0
M2 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=3990 $Y=660 $dt=0
M3 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=6470 $Y=660 $dt=0
M4 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=8950 $Y=660 $dt=0
M5 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=4.312e-13 AS=2.376e-13 PD=2.74e-06 PS=1.42e-06 $X=11430 $Y=660 $dt=0
M6 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.5505e-13 AS=6.312e-13 PD=1.855e-06 PS=3.59e-06 $X=620 $Y=2505 $dt=1
M7 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.5505e-13 AS=3.5505e-13 PD=1.855e-06 PS=1.855e-06 $X=3090 $Y=2505 $dt=1
M8 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.5505e-13 AS=3.5505e-13 PD=1.855e-06 PS=1.855e-06 $X=5560 $Y=2505 $dt=1
M9 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.5505e-13 AS=3.5505e-13 PD=1.855e-06 PS=1.855e-06 $X=8030 $Y=2505 $dt=1
M10 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.84638e-13 AS=3.5505e-13 PD=1.9e-06 PS=1.855e-06 $X=10500 $Y=2505 $dt=1
M11 5 4 vdd3i! vdd3i! pe3i L=3e-07 W=1.315e-06 AD=7.56575e-13 AS=3.84638e-13 PD=3.91e-06 PS=1.9e-06 $X=13015 $Y=2505 $dt=1
.ends DECAP25JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP15JI3V                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP15JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=8
M0 gnd3i! 5 4 gnd3i! ne3i L=3.5e-07 W=8.8e-07 AD=2.42e-13 AS=4.224e-13 PD=1.43e-06 PS=2.72e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.71e-06 W=8.8e-07 AD=2.42e-13 AS=2.42e-13 PD=1.43e-06 PS=1.43e-06 $X=1520 $Y=660 $dt=0
M2 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.71e-06 W=8.8e-07 AD=2.376e-13 AS=2.42e-13 PD=1.42e-06 PS=1.43e-06 $X=3780 $Y=660 $dt=0
M3 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.71e-06 W=8.8e-07 AD=6.046e-13 AS=2.376e-13 PD=3.5e-06 PS=1.42e-06 $X=6030 $Y=660 $dt=0
M4 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.7e-06 W=1.315e-06 AD=3.5505e-13 AS=8.308e-13 PD=1.855e-06 PS=4.37e-06 $X=660 $Y=2505 $dt=1
M5 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.7e-06 W=1.315e-06 AD=3.5505e-13 AS=3.5505e-13 PD=1.855e-06 PS=1.855e-06 $X=2900 $Y=2505 $dt=1
M6 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.7e-06 W=1.315e-06 AD=3.78063e-13 AS=3.5505e-13 PD=1.89e-06 PS=1.855e-06 $X=5140 $Y=2505 $dt=1
M7 5 4 vdd3i! vdd3i! pe3i L=3e-07 W=1.315e-06 AD=7.56575e-13 AS=3.78063e-13 PD=3.91e-06 PS=1.89e-06 $X=7415 $Y=2505 $dt=1
.ends DECAP15JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP7JI3V                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP7JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=4
M0 gnd3i! 5 4 gnd3i! ne3i L=3.5e-07 W=8.8e-07 AD=2.376e-13 AS=4.224e-13 PD=1.42e-06 PS=2.72e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.75e-06 W=8.8e-07 AD=6.046e-13 AS=2.376e-13 PD=3.5e-06 PS=1.42e-06 $X=1510 $Y=660 $dt=0
M2 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.71e-06 W=1.315e-06 AD=3.87925e-13 AS=8.308e-13 PD=1.905e-06 PS=4.37e-06 $X=660 $Y=2505 $dt=1
M3 5 4 vdd3i! vdd3i! pe3i L=3e-07 W=1.315e-06 AD=7.237e-13 AS=3.87925e-13 PD=3.86e-06 PS=1.905e-06 $X=2960 $Y=2505 $dt=1
.ends DECAP7JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP5JI3V                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP5JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=2
M0 gnd3i! 5 4 gnd3i! ne3i L=1.48e-06 W=8.3e-07 AD=5.786e-13 AS=4.568e-13 PD=3.4e-06 PS=2.82e-06 $X=660 $Y=660 $dt=0
M1 5 4 vdd3i! vdd3i! pe3i L=1.46e-06 W=1.36e-06 AD=7.564e-13 AS=8.542e-13 PD=3.9e-06 PS=4.46e-06 $X=660 $Y=2460 $dt=1
.ends DECAP5JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP10JI3V                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP10JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=6
M0 gnd3i! 5 4 gnd3i! ne3i L=3.5e-07 W=8.8e-07 AD=2.376e-13 AS=4.224e-13 PD=1.42e-06 PS=2.72e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.445e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=1510 $Y=660 $dt=0
M2 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.445e-06 W=8.8e-07 AD=6.046e-13 AS=2.376e-13 PD=3.5e-06 PS=1.42e-06 $X=3495 $Y=660 $dt=0
M3 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.425e-06 W=1.315e-06 AD=3.5505e-13 AS=8.308e-13 PD=1.855e-06 PS=4.37e-06 $X=660 $Y=2505 $dt=1
M4 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.425e-06 W=1.315e-06 AD=3.71488e-13 AS=3.5505e-13 PD=1.88e-06 PS=1.855e-06 $X=2625 $Y=2505 $dt=1
M5 5 4 vdd3i! vdd3i! pe3i L=3e-07 W=1.315e-06 AD=7.56575e-13 AS=3.71488e-13 PD=3.91e-06 PS=1.88e-06 $X=4615 $Y=2505 $dt=1
.ends DECAP10JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: aska_dig                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt aska_dig 1 2 enable DAC<0> pulse_active DAC<1> DAC<2> DAC<4> DAC<3> down_switches<4>
+ down_switches<1> down_switches<2> down_switches<3> SPI_CS down_switches<5> down_switches<6> SPI_Clk down_switches<7> down_switches<9> down_switches<8>
+ down_switches<10> down_switches<0> down_switches<11> down_switches<14> down_switches<12> DAC<5> clk down_switches<13> up_switches<0> down_switches<15>
+ reset_l up_switches<9> up_switches<6> up_switches<8> porborn up_switches<3> up_switches<2> down_switches<17> down_switches<16> up_switches<1>
+ up_switches<4> up_switches<10> SPI_MOSI down_switches<20> up_switches<7> down_switches<18> down_switches<19> up_switches<5> up_switches<12> up_switches<11>
+ IC_addr<1> down_switches<21> up_switches<13> down_switches<22> IC_addr<0> up_switches<14> up_switches<15> down_switches<23> down_switches<24> up_switches<22>
+ up_switches<16> down_switches<25> up_switches<17> up_switches<18> up_switches<19> down_switches<26> up_switches<21> down_switches<27> up_switches<20> down_switches<28>
+ up_switches<23> up_switches<26> up_switches<25> down_switches<31> up_switches<24> up_switches<27> up_switches<28> down_switches<30> down_switches<29> up_switches<29>
+ up_switches<30> up_switches<31>
** N=1434 EP=82 FDC=26952
X8325 1 2 162 1172 170 EN2JI3VX0 $T=40320 185920 1 0 $X=39890 $Y=180800
X8326 1 2 173 706 754 EN2JI3VX0 $T=45920 185920 1 0 $X=45490 $Y=180800
X8327 1 2 555 546 922 EN2JI3VX0 $T=306880 212800 1 180 $X=300850 $Y=212160
X8328 1 2 1140 615 1316 621 NO3JI3VX1 $T=347760 24640 1 180 $X=343970 $Y=24000
X8329 1 2 537 111 1130 NA2JI3VX2 $T=307440 105280 0 0 $X=307010 $Y=104640
X8330 1 2 1123 589 1293 585 NO22JI3VX1 $T=328160 168000 0 180 $X=323250 $Y=162880
X8331 1 2 966 662 1161 1365 NO22JI3VX1 $T=397040 141120 1 180 $X=392130 $Y=140480
X8332 1 2 590 1135 116 593 DFRRQJI3VX2 $T=342720 212800 0 180 $X=326050 $Y=207680
X8333 1 2 1366 DAC<0> BUJI3VX8 $T=50960 33600 1 0 $X=50530 $Y=28480
X8334 1 2 1367 DAC<4> BUJI3VX8 $T=67200 33600 1 0 $X=66770 $Y=28480
X8335 1 2 231 258 BUJI3VX8 $T=91280 141120 1 0 $X=90850 $Y=136000
X8336 1 2 231 257 BUJI3VX8 $T=103600 168000 1 0 $X=103170 $Y=162880
X8337 1 2 267 84 BUJI3VX8 $T=126560 203840 0 180 $X=117730 $Y=198720
X8338 1 2 267 92 BUJI3VX8 $T=175280 114240 0 0 $X=174850 $Y=113600
X8339 1 2 357 DAC<5> BUJI3VX8 $T=176400 24640 1 0 $X=175970 $Y=19520
X8340 1 2 267 98 BUJI3VX8 $T=218400 203840 0 0 $X=217970 $Y=203200
X8341 1 2 267 102 BUJI3VX8 $T=314720 194880 1 0 $X=314290 $Y=189760
X8342 1 2 442 1335 98 515 DFRRQJI3VX4 $T=297360 176960 1 180 $X=279010 $Y=176320
X8343 1 2 590 619 116 622 DFRRQJI3VX4 $T=334880 203840 1 0 $X=334450 $Y=198720
X8344 1 2 105 955 102 954 DFRRQJI3VX4 $T=379120 185920 1 180 $X=360770 $Y=185280
X8345 1 2 105 649 102 661 DFRRQJI3VX4 $T=371840 168000 0 0 $X=371410 $Y=167360
X8346 1 2 105 969 102 1159 DFRRQJI3VX4 $T=407680 168000 1 180 $X=389330 $Y=167360
X8347 1 2 105 974 102 670 DFRRQJI3VX4 $T=413840 123200 1 180 $X=395490 $Y=122560
X8348 1 2 105 1314 102 693 DFRRQJI3VX4 $T=416080 123200 0 180 $X=397730 $Y=118080
X8349 1 2 742 775 BUJI3VX1 $T=36960 176960 0 0 $X=36530 $Y=176320
X8350 1 2 SPI_Clk 496 BUJI3VX1 $T=120400 96320 0 0 $X=119970 $Y=95680
X8351 1 2 clk 611 BUJI3VX1 $T=186480 159040 0 0 $X=186050 $Y=158400
X8352 1 2 123 109 BUJI3VX1 $T=207200 87360 1 0 $X=206770 $Y=82240
X8353 1 2 417 123 BUJI3VX1 $T=207200 212800 0 0 $X=206770 $Y=212160
X8354 1 2 525 126 BUJI3VX1 $T=208320 194880 1 0 $X=207890 $Y=189760
X8355 1 2 1076 861 BUJI3VX1 $T=211120 194880 1 0 $X=210690 $Y=189760
X8356 1 2 496 742 BUJI3VX1 $T=270480 203840 0 180 $X=267250 $Y=198720
X8357 1 2 611 494 BUJI3VX1 $T=339360 185920 0 180 $X=336130 $Y=180800
X8358 1 2 521 690 BUJI3VX1 $T=403760 105280 0 0 $X=403330 $Y=104640
X8359 1 2 718 127 408 319 NO3I2JI3VX1 $T=209440 185920 1 180 $X=205090 $Y=185280
X8360 1 2 97 859 133 1116 NO3I2JI3VX1 $T=220080 176960 0 0 $X=219650 $Y=176320
X8361 1 2 272 278 1019 260 794 FAJI3VX1 $T=112000 168000 1 0 $X=111570 $Y=162880
X8362 1 2 804 794 1017 1011 263 FAJI3VX1 $T=129360 159040 1 180 $X=114370 $Y=158400
X8363 1 2 803 263 296 808 269 FAJI3VX1 $T=133840 150080 0 180 $X=118850 $Y=144960
X8364 1 2 1014 281 1018 806 278 FAJI3VX1 $T=123200 185920 0 0 $X=122770 $Y=185280
X8365 1 2 1024 282 798 821 274 FAJI3VX1 $T=137760 212800 0 180 $X=122770 $Y=207680
X8366 1 2 1028 274 1016 264 281 FAJI3VX1 $T=141120 203840 0 180 $X=126130 $Y=198720
X8367 1 2 308 1213 321 808 317 FAJI3VX1 $T=150640 150080 0 180 $X=135650 $Y=144960
X8368 1 2 1219 977 302 1011 1213 FAJI3VX1 $T=150640 150080 1 180 $X=135650 $Y=149440
X8369 1 2 814 298 291 260 977 FAJI3VX1 $T=151200 168000 0 180 $X=136210 $Y=162880
X8370 1 2 292 301 118 806 298 FAJI3VX1 $T=137760 185920 0 0 $X=137330 $Y=185280
X8371 1 2 1029 816 1217 821 305 FAJI3VX1 $T=140560 212800 0 0 $X=140130 $Y=212160
X8372 1 2 1040 305 1030 264 301 FAJI3VX1 $T=155680 203840 0 180 $X=140690 $Y=198720
X8373 1 2 315 824 820 1368 328 FAJI3VX1 $T=148400 114240 0 0 $X=147970 $Y=113600
X8374 1 2 827 269 309 307 345 FAJI3VX1 $T=164640 141120 1 180 $X=149650 $Y=140480
X8375 1 2 330 317 820 307 346 FAJI3VX1 $T=166320 150080 1 180 $X=151330 $Y=149440
X8376 1 2 833 328 333 324 1051 FAJI3VX1 $T=175840 123200 0 180 $X=160850 $Y=118080
X8377 1 2 1320 345 335 329 354 FAJI3VX1 $T=180320 141120 0 180 $X=165330 $Y=136000
X8378 1 2 830 346 333 329 359 FAJI3VX1 $T=181440 150080 1 180 $X=166450 $Y=149440
X8379 1 2 844 368 849 OR2JI3VX0 $T=183680 194880 0 0 $X=183250 $Y=194240
X8380 1 2 425 220 129 OR2JI3VX0 $T=208880 168000 0 0 $X=208450 $Y=167360
X8381 1 2 448 1103 1099 OR2JI3VX0 $T=240800 168000 0 0 $X=240370 $Y=167360
X8382 1 2 544 220 1286 OR2JI3VX0 $T=303520 168000 1 0 $X=303090 $Y=162880
X8383 1 2 447 609 695 OR2JI3VX0 $T=388080 159040 1 0 $X=387650 $Y=153920
X8384 1 2 163 1369 160 165 NA3I1JI3VX1 $T=36960 150080 0 0 $X=36530 $Y=149440
X8385 1 2 767 1359 995 996 NA3I1JI3VX1 $T=61040 176960 0 0 $X=60610 $Y=176320
X8386 1 2 765 539 202 1370 NA3I1JI3VX1 $T=64400 168000 1 0 $X=63970 $Y=162880
X8387 1 2 764 765 766 179 NA3I1JI3VX1 $T=68880 159040 1 180 $X=64530 $Y=158400
X8388 1 2 593 556 576 613 NA3I1JI3VX1 $T=329280 212800 1 180 $X=324930 $Y=212160
X8389 1 2 939 1298 582 935 NA3I1JI3VX1 $T=337680 168000 0 180 $X=333330 $Y=162880
X8390 1 2 661 1371 683 1159 NA3I1JI3VX1 $T=386960 168000 1 0 $X=386530 $Y=162880
X8391 1 2 670 1372 693 681 NA3I1JI3VX1 $T=395920 114240 1 180 $X=391570 $Y=113600
X8392 1 2 690 972 1166 693 NA3I1JI3VX1 $T=401520 114240 1 0 $X=401090 $Y=109120
X8393 1 2 231 248 DLY2JI3VX1 $T=77840 212800 0 0 $X=77410 $Y=212160
X8394 1 2 152 163 1171 150 NA3JI3VX0 $T=40320 168000 0 180 $X=37090 $Y=162880
X8395 1 2 1373 178 757 110 NA3JI3VX0 $T=57120 159040 1 180 $X=53890 $Y=158400
X8396 1 2 1374 195 186 194 NA3JI3VX0 $T=58240 150080 0 0 $X=57810 $Y=149440
X8397 1 2 152 87 210 212 NA3JI3VX0 $T=67760 185920 0 0 $X=67330 $Y=185280
X8398 1 2 212 199 772 203 NA3JI3VX0 $T=75600 194880 0 180 $X=72370 $Y=189760
X8399 1 2 1020 807 1025 300 NA3JI3VX0 $T=133280 123200 1 0 $X=132850 $Y=118080
X8400 1 2 295 293 1375 90 NA3JI3VX0 $T=141120 114240 0 0 $X=140690 $Y=113600
X8401 1 2 120 823 119 1044 NA3JI3VX0 $T=154560 105280 0 0 $X=154130 $Y=104640
X8402 1 2 382 358 384 127 NA3JI3VX0 $T=194320 176960 0 180 $X=191090 $Y=171840
X8403 1 2 1069 1067 385 1236 NA3JI3VX0 $T=194320 185920 1 180 $X=191090 $Y=185280
X8404 1 2 1068 401 852 1073 NA3JI3VX0 $T=196560 203840 1 0 $X=196130 $Y=198720
X8405 1 2 1170 433 883 134 NA3JI3VX0 $T=240800 185920 1 180 $X=237570 $Y=185280
X8406 1 2 1376 469 464 467 NA3JI3VX0 $T=250320 159040 0 0 $X=249890 $Y=158400
X8407 1 2 127 485 904 906 NA3JI3VX0 $T=271040 185920 1 0 $X=270610 $Y=180800
X8408 1 2 160 178 1176 983 ON21JI3VX1 $T=36960 159040 0 180 $X=33170 $Y=153920
X8409 1 2 152 1176 1177 756 ON21JI3VX1 $T=38640 159040 1 0 $X=38210 $Y=153920
X8410 1 2 1189 198 1317 761 ON21JI3VX1 $T=62720 168000 1 180 $X=58930 $Y=167360
X8411 1 2 210 219 1318 87 ON21JI3VX1 $T=72800 185920 0 0 $X=72370 $Y=185280
X8412 1 2 361 1377 1232 847 ON21JI3VX1 $T=180880 176960 0 0 $X=180450 $Y=176320
X8413 1 2 1378 358 1345 846 ON21JI3VX1 $T=191520 168000 1 180 $X=187730 $Y=167360
X8414 1 2 1070 1065 851 385 ON21JI3VX1 $T=194320 185920 1 0 $X=193890 $Y=180800
X8415 1 2 129 857 1324 1246 ON21JI3VX1 $T=202720 168000 1 0 $X=202290 $Y=162880
X8416 1 2 220 421 1379 1244 ON21JI3VX1 $T=209440 176960 0 180 $X=205650 $Y=171840
X8417 1 2 1080 130 423 856 ON21JI3VX1 $T=210560 185920 0 0 $X=210130 $Y=185280
X8418 1 2 1086 1347 876 1250 ON21JI3VX1 $T=218960 203840 1 0 $X=218530 $Y=198720
X8419 1 2 883 1100 1252 433 ON21JI3VX1 $T=237440 185920 1 180 $X=233650 $Y=185280
X8420 1 2 886 1093 1380 1099 ON21JI3VX1 $T=241920 159040 0 0 $X=241490 $Y=158400
X8421 1 2 1098 467 1101 889 ON21JI3VX1 $T=249760 168000 0 180 $X=245970 $Y=162880
X8422 1 2 466 885 894 1105 ON21JI3VX1 $T=250320 168000 0 0 $X=249890 $Y=167360
X8423 1 2 447 897 584 1334 ON21JI3VX1 $T=258160 33600 0 0 $X=257730 $Y=32960
X8424 1 2 220 1116 1381 1244 ON21JI3VX1 $T=264880 176960 0 0 $X=264450 $Y=176320
X8425 1 2 1382 485 1335 511 ON21JI3VX1 $T=285600 185920 0 180 $X=281810 $Y=180800
X8426 1 2 447 914 605 907 ON21JI3VX1 $T=283920 33600 0 0 $X=283490 $Y=32960
X8427 1 2 447 528 917 913 ON21JI3VX1 $T=285040 24640 0 0 $X=284610 $Y=24000
X8428 1 2 928 1383 557 1289 ON21JI3VX1 $T=317520 168000 1 180 $X=313730 $Y=167360
X8429 1 2 447 138 944 1303 ON21JI3VX1 $T=337680 33600 0 0 $X=337250 $Y=32960
X8430 1 2 447 1384 953 951 ON21JI3VX1 $T=348880 42560 1 0 $X=348450 $Y=37440
X8431 1 2 1144 948 955 142 ON21JI3VX1 $T=360080 185920 1 0 $X=359650 $Y=180800
X8432 1 2 447 1356 1148 1355 ON21JI3VX1 $T=371280 33600 1 180 $X=367490 $Y=32960
X8433 1 2 447 1156 658 1339 ON21JI3VX1 $T=376880 24640 0 0 $X=376450 $Y=24000
X8434 1 2 1371 981 649 665 ON21JI3VX1 $T=384720 168000 0 180 $X=380930 $Y=162880
X8435 1 2 1159 1358 1385 685 ON21JI3VX1 $T=390880 159040 1 180 $X=387090 $Y=158400
X8436 1 2 682 1365 960 680 ON21JI3VX1 $T=391440 141120 1 180 $X=387650 $Y=140480
X8437 1 2 1386 676 1357 670 ON21JI3VX1 $T=388640 114240 0 0 $X=388210 $Y=113600
X8438 1 2 683 1358 1165 695 ON21JI3VX1 $T=392000 159040 1 0 $X=391570 $Y=153920
X8439 1 2 1372 145 974 1357 ON21JI3VX1 $T=397600 114240 0 0 $X=397170 $Y=113600
X8440 1 2 693 145 1314 972 ON21JI3VX1 $T=403760 114240 0 0 $X=403330 $Y=113600
X8441 1 2 998 996 767 198 OA21JI3VX1 $T=69440 176960 1 180 $X=64530 $Y=176320
X8442 1 2 546 566 577 1131 OA21JI3VX1 $T=316400 212800 0 0 $X=315970 $Y=212160
X8443 1 2 231 244 BUJI3VX3 $T=110320 203840 1 0 $X=109890 $Y=198720
X8444 1 2 231 247 BUJI3VX3 $T=113680 212800 1 0 $X=113250 $Y=207680
X8445 1 2 231 1013 BUJI3VX3 $T=119280 212800 1 0 $X=118850 $Y=207680
X8446 1 2 231 285 BUJI3VX3 $T=136640 176960 1 0 $X=136210 $Y=171840
X8447 1 2 231 287 BUJI3VX3 $T=137200 168000 0 0 $X=136770 $Y=167360
X8448 1 2 231 280 BUJI3VX3 $T=137760 185920 1 0 $X=137330 $Y=180800
X8449 1 2 231 406 BUJI3VX3 $T=189280 159040 0 0 $X=188850 $Y=158400
X8450 1 2 397 up_switches<0> BUJI3VX3 $T=203840 24640 1 0 $X=203410 $Y=19520
X8451 1 2 415 up_switches<9> BUJI3VX3 $T=208880 24640 1 0 $X=208450 $Y=19520
X8452 1 2 422 up_switches<8> BUJI3VX3 $T=213360 24640 1 0 $X=212930 $Y=19520
X8453 1 2 405 up_switches<6> BUJI3VX3 $T=213360 24640 0 0 $X=212930 $Y=24000
X8454 1 2 429 up_switches<3> BUJI3VX3 $T=221200 24640 1 180 $X=216850 $Y=24000
X8455 1 2 221 up_switches<2> BUJI3VX3 $T=217840 24640 1 0 $X=217410 $Y=19520
X8456 1 2 231 871 BUJI3VX3 $T=220640 168000 1 0 $X=220210 $Y=162880
X8457 1 2 432 468 BUJI3VX3 $T=220640 194880 1 0 $X=220210 $Y=189760
X8458 1 2 231 868 BUJI3VX3 $T=234640 150080 0 180 $X=230290 $Y=144960
X8459 1 2 468 525 BUJI3VX3 $T=233520 176960 1 0 $X=233090 $Y=171840
X8460 1 2 222 up_switches<1> BUJI3VX3 $T=240800 24640 1 0 $X=240370 $Y=19520
X8461 1 2 451 up_switches<4> BUJI3VX3 $T=245840 24640 1 0 $X=245410 $Y=19520
X8462 1 2 460 up_switches<10> BUJI3VX3 $T=253120 24640 1 0 $X=252690 $Y=19520
X8463 1 2 231 454 BUJI3VX3 $T=255360 123200 0 0 $X=254930 $Y=122560
X8464 1 2 409 up_switches<7> BUJI3VX3 $T=258720 24640 1 0 $X=258290 $Y=19520
X8465 1 2 484 up_switches<5> BUJI3VX3 $T=264880 24640 1 0 $X=264450 $Y=19520
X8466 1 2 499 up_switches<12> BUJI3VX3 $T=271600 24640 1 0 $X=271170 $Y=19520
X8467 1 2 353 up_switches<11> BUJI3VX3 $T=277200 24640 1 0 $X=276770 $Y=19520
X8468 1 2 419 up_switches<13> BUJI3VX3 $T=282240 24640 1 0 $X=281810 $Y=19520
X8469 1 2 746 991 174 172 1178 AN211JI3VX1 $T=45360 168000 0 0 $X=44930 $Y=167360
X8470 1 2 186 764 1373 220 197 AN211JI3VX1 $T=64400 159040 1 180 $X=59490 $Y=158400
X8471 1 2 1387 343 853 1070 1388 AN211JI3VX1 $T=193200 176960 0 0 $X=192770 $Y=176320
X8472 1 2 423 131 408 1088 425 AN211JI3VX1 $T=217280 185920 0 180 $X=212370 $Y=180800
X8473 1 2 617 612 1289 618 140 AN211JI3VX1 $T=343280 168000 0 180 $X=338370 $Y=162880
X8474 1 2 231 255 BUJI3VX16 $T=110320 203840 0 180 $X=93650 $Y=198720
X8475 1 2 826 380 BUJI3VX16 $T=159600 203840 1 0 $X=159170 $Y=198720
X8476 1 2 231 387 BUJI3VX16 $T=210000 123200 1 0 $X=209570 $Y=118080
X8477 1 2 231 306 BUJI3VX16 $T=239680 132160 0 180 $X=223010 $Y=127040
X8478 1 2 153 165 BUJI3VX0 $T=44240 150080 0 0 $X=43810 $Y=149440
X8479 1 2 168 990 BUJI3VX0 $T=44240 159040 1 0 $X=43810 $Y=153920
X8480 1 2 173 993 BUJI3VX0 $T=54880 194880 1 0 $X=54450 $Y=189760
X8481 1 2 708 994 BUJI3VX0 $T=62720 185920 1 0 $X=62290 $Y=180800
X8482 1 2 819 1218 BUJI3VX0 $T=151200 114240 1 0 $X=150770 $Y=109120
X8483 1 2 825 1361 BUJI3VX0 $T=161840 114240 1 0 $X=161410 $Y=109120
X8484 1 2 823 327 BUJI3VX0 $T=162400 96320 1 0 $X=161970 $Y=91200
X8485 1 2 316 340 BUJI3VX0 $T=165760 212800 1 0 $X=165330 $Y=207680
X8486 1 2 828 1047 BUJI3VX0 $T=190400 105280 0 0 $X=189970 $Y=104640
X8487 1 2 126 1076 BUJI3VX0 $T=204960 194880 0 0 $X=204530 $Y=194240
X8488 1 2 861 431 BUJI3VX0 $T=207760 194880 0 0 $X=207330 $Y=194240
X8489 1 2 864 1327 BUJI3VX0 $T=213920 194880 1 0 $X=213490 $Y=189760
X8490 1 2 1327 865 BUJI3VX0 $T=215040 203840 1 0 $X=214610 $Y=198720
X8491 1 2 870 864 BUJI3VX0 $T=215600 203840 0 0 $X=215170 $Y=203200
X8492 1 2 porborn 870 BUJI3VX0 $T=218400 212800 0 0 $X=217970 $Y=212160
X8493 1 2 1102 432 BUJI3VX0 $T=231840 203840 1 0 $X=231410 $Y=198720
X8494 1 2 440 134 BUJI3VX0 $T=238000 176960 1 0 $X=237570 $Y=171840
X8495 1 2 882 887 BUJI3VX0 $T=241920 203840 0 0 $X=241490 $Y=203200
X8496 1 2 892 891 BUJI3VX0 $T=244720 185920 0 0 $X=244290 $Y=185280
X8497 1 2 887 1102 BUJI3VX0 $T=244720 212800 1 0 $X=244290 $Y=207680
X8498 1 2 SPI_MOSI 1269 BUJI3VX0 $T=260400 212800 0 0 $X=259970 $Y=212160
X8499 1 2 900 882 BUJI3VX0 $T=264320 212800 1 0 $X=263890 $Y=207680
X8500 1 2 529 536 BUJI3VX0 $T=288960 185920 0 0 $X=288530 $Y=185280
X8501 1 2 541 919 BUJI3VX0 $T=295680 194880 1 0 $X=295250 $Y=189760
X8502 1 2 922 923 BUJI3VX0 $T=302400 203840 0 0 $X=301970 $Y=203200
X8503 1 2 559 577 BUJI3VX0 $T=320880 212800 0 0 $X=320450 $Y=212160
X8504 1 2 730 1389 BUJI3VX0 $T=349440 212800 0 0 $X=349010 $Y=212160
X8505 1 2 1172 986 162 NA2I1JI3VX1 $T=47600 176960 1 180 $X=43810 $Y=176320
X8506 1 2 706 1172 173 NA2I1JI3VX1 $T=50960 176960 1 180 $X=47170 $Y=176320
X8507 1 2 182 194 756 NA2I1JI3VX1 $T=57680 150080 1 180 $X=53890 $Y=149440
X8508 1 2 756 186 182 NA2I1JI3VX1 $T=54320 159040 1 0 $X=53890 $Y=153920
X8509 1 2 1390 763 994 NA2I1JI3VX1 $T=59360 185920 0 0 $X=58930 $Y=185280
X8510 1 2 819 1035 302 NA2I1JI3VX1 $T=142240 132160 1 0 $X=141810 $Y=127040
X8511 1 2 303 1216 1035 NA2I1JI3VX1 $T=150080 123200 1 180 $X=146290 $Y=122560
X8512 1 2 320 1391 91 NA2I1JI3VX1 $T=160720 132160 0 180 $X=156930 $Y=127040
X8513 1 2 828 91 321 NA2I1JI3VX1 $T=162960 123200 1 180 $X=159170 $Y=122560
X8514 1 2 1058 840 361 NA2I1JI3VX1 $T=176960 185920 1 0 $X=176530 $Y=180800
X8515 1 2 364 385 1071 NA2I1JI3VX1 $T=194880 194880 1 0 $X=194450 $Y=189760
X8516 1 2 1071 1073 395 NA2I1JI3VX1 $T=196000 212800 0 0 $X=195570 $Y=212160
X8517 1 2 1071 391 364 NA2I1JI3VX1 $T=201600 194880 0 180 $X=197810 $Y=189760
X8518 1 2 395 852 1071 NA2I1JI3VX1 $T=199360 203840 1 0 $X=198930 $Y=198720
X8519 1 2 407 399 426 NA2I1JI3VX1 $T=204960 176960 0 180 $X=201170 $Y=171840
X8520 1 2 97 420 1392 NA2I1JI3VX1 $T=214480 176960 0 180 $X=210690 $Y=171840
X8521 1 2 859 720 133 NA2I1JI3VX1 $T=219520 168000 0 0 $X=219090 $Y=167360
X8522 1 2 720 544 97 NA2I1JI3VX1 $T=223440 176960 0 180 $X=219650 $Y=171840
X8523 1 2 1263 1257 891 NA2I1JI3VX1 $T=250320 194880 0 180 $X=246530 $Y=189760
X8524 1 2 505 1393 487 NA2I1JI3VX1 $T=268240 168000 0 180 $X=264450 $Y=162880
X8525 1 2 905 498 495 NA2I1JI3VX1 $T=272720 168000 1 180 $X=268930 $Y=167360
X8526 1 2 515 495 518 NA2I1JI3VX1 $T=276640 168000 1 180 $X=272850 $Y=167360
X8527 1 2 909 487 506 NA2I1JI3VX1 $T=276640 176960 1 180 $X=272850 $Y=176320
X8528 1 2 610 575 591 NA2I1JI3VX1 $T=322560 176960 0 180 $X=318770 $Y=171840
X8529 1 2 591 586 610 NA2I1JI3VX1 $T=328160 176960 1 0 $X=327730 $Y=171840
X8530 1 2 601 946 600 NA2I1JI3VX1 $T=334320 176960 0 0 $X=333890 $Y=176320
X8531 1 2 703 984 DLY1JI3VX1 $T=28560 141120 1 0 $X=28130 $Y=136000
X8532 1 2 146 741 DLY1JI3VX1 $T=29680 114240 0 0 $X=29250 $Y=113600
X8533 1 2 704 740 DLY1JI3VX1 $T=29680 123200 1 0 $X=29250 $Y=118080
X8534 1 2 158 743 DLY1JI3VX1 $T=34160 141120 1 0 $X=33730 $Y=136000
X8535 1 2 159 744 DLY1JI3VX1 $T=34160 141120 0 0 $X=33730 $Y=140480
X8536 1 2 187 1179 DLY1JI3VX1 $T=44240 33600 0 0 $X=43810 $Y=32960
X8537 1 2 987 1181 DLY1JI3VX1 $T=47040 123200 0 0 $X=46610 $Y=122560
X8538 1 2 705 1183 DLY1JI3VX1 $T=49840 33600 0 0 $X=49410 $Y=32960
X8539 1 2 185 1187 DLY1JI3VX1 $T=56000 33600 0 0 $X=55570 $Y=32960
X8540 1 2 1003 1190 DLY1JI3VX1 $T=61600 33600 0 0 $X=61170 $Y=32960
X8541 1 2 1193 1000 DLY1JI3VX1 $T=65520 150080 0 0 $X=65090 $Y=149440
X8542 1 2 709 1192 DLY1JI3VX1 $T=67200 33600 0 0 $X=66770 $Y=32960
X8543 1 2 1001 1002 DLY1JI3VX1 $T=69440 69440 1 0 $X=69010 $Y=64320
X8544 1 2 768 1194 DLY1JI3VX1 $T=72240 141120 0 0 $X=71810 $Y=140480
X8545 1 2 218 774 DLY1JI3VX1 $T=72800 33600 0 0 $X=72370 $Y=32960
X8546 1 2 710 1196 DLY1JI3VX1 $T=78400 33600 0 0 $X=77970 $Y=32960
X8547 1 2 1198 229 DLY1JI3VX1 $T=84560 185920 0 0 $X=84130 $Y=185280
X8548 1 2 711 785 DLY1JI3VX1 $T=85120 87360 1 0 $X=84690 $Y=82240
X8549 1 2 225 781 DLY1JI3VX1 $T=85120 203840 1 0 $X=84690 $Y=198720
X8550 1 2 788 234 DLY1JI3VX1 $T=87360 168000 1 0 $X=86930 $Y=162880
X8551 1 2 780 235 DLY1JI3VX1 $T=87360 168000 0 0 $X=86930 $Y=167360
X8552 1 2 712 1168 DLY1JI3VX1 $T=89040 150080 1 0 $X=88610 $Y=144960
X8553 1 2 782 1197 DLY1JI3VX1 $T=95200 203840 1 180 $X=89170 $Y=203200
X8554 1 2 246 1201 DLY1JI3VX1 $T=103040 203840 0 0 $X=102610 $Y=203200
X8555 1 2 1199 1008 DLY1JI3VX1 $T=103600 69440 0 0 $X=103170 $Y=68800
X8556 1 2 1202 1010 DLY1JI3VX1 $T=108640 159040 0 0 $X=108210 $Y=158400
X8557 1 2 256 1012 DLY1JI3VX1 $T=113680 150080 1 0 $X=113250 $Y=144960
X8558 1 2 789 795 DLY1JI3VX1 $T=113680 168000 0 0 $X=113250 $Y=167360
X8559 1 2 792 797 DLY1JI3VX1 $T=117040 33600 1 0 $X=116610 $Y=28480
X8560 1 2 790 1022 DLY1JI3VX1 $T=129360 42560 1 0 $X=128930 $Y=37440
X8561 1 2 1204 1023 DLY1JI3VX1 $T=132160 185920 1 0 $X=131730 $Y=180800
X8562 1 2 1009 1209 DLY1JI3VX1 $T=134960 42560 1 0 $X=134530 $Y=37440
X8563 1 2 1203 1027 DLY1JI3VX1 $T=134960 132160 0 0 $X=134530 $Y=131520
X8564 1 2 800 811 DLY1JI3VX1 $T=136080 69440 0 0 $X=135650 $Y=68800
X8565 1 2 791 1031 DLY1JI3VX1 $T=140560 42560 1 0 $X=140130 $Y=37440
X8566 1 2 715 1215 DLY1JI3VX1 $T=140560 132160 0 0 $X=140130 $Y=131520
X8567 1 2 802 1220 DLY1JI3VX1 $T=146160 42560 1 0 $X=145730 $Y=37440
X8568 1 2 1034 1039 DLY1JI3VX1 $T=146160 60480 1 0 $X=145730 $Y=55360
X8569 1 2 1360 88 DLY1JI3VX1 $T=146160 132160 0 0 $X=145730 $Y=131520
X8570 1 2 1032 1041 DLY1JI3VX1 $T=151760 60480 1 0 $X=151330 $Y=55360
X8571 1 2 813 1222 DLY1JI3VX1 $T=152880 42560 1 0 $X=152450 $Y=37440
X8572 1 2 1045 1225 DLY1JI3VX1 $T=157360 60480 1 0 $X=156930 $Y=55360
X8573 1 2 1048 1226 DLY1JI3VX1 $T=158480 42560 1 0 $X=158050 $Y=37440
X8574 1 2 1052 1054 DLY1JI3VX1 $T=167440 114240 1 0 $X=167010 $Y=109120
X8575 1 2 1059 1227 DLY1JI3VX1 $T=169120 33600 0 0 $X=168690 $Y=32960
X8576 1 2 1228 1229 DLY1JI3VX1 $T=174720 33600 0 0 $X=174290 $Y=32960
X8577 1 2 1056 1323 DLY1JI3VX1 $T=174720 132160 1 0 $X=174290 $Y=127040
X8578 1 2 375 1231 DLY1JI3VX1 $T=177520 96320 0 0 $X=177090 $Y=95680
X8579 1 2 836 1233 DLY1JI3VX1 $T=179200 42560 1 0 $X=178770 $Y=37440
X8580 1 2 1082 1235 DLY1JI3VX1 $T=186480 141120 1 0 $X=186050 $Y=136000
X8581 1 2 1072 1237 DLY1JI3VX1 $T=187600 42560 1 0 $X=187170 $Y=37440
X8582 1 2 717 1239 DLY1JI3VX1 $T=190960 105280 1 0 $X=190530 $Y=100160
X8583 1 2 383 1240 DLY1JI3VX1 $T=192080 33600 0 0 $X=191650 $Y=32960
X8584 1 2 1083 1241 DLY1JI3VX1 $T=192080 132160 0 0 $X=191650 $Y=131520
X8585 1 2 1066 1242 DLY1JI3VX1 $T=193200 105280 0 0 $X=192770 $Y=104640
X8586 1 2 394 403 DLY1JI3VX1 $T=197680 123200 1 0 $X=197250 $Y=118080
X8587 1 2 1234 1075 DLY1JI3VX1 $T=197680 132160 0 0 $X=197250 $Y=131520
X8588 1 2 SPI_CS 826 DLY1JI3VX1 $T=201600 212800 0 0 $X=201170 $Y=212160
X8589 1 2 719 424 DLY1JI3VX1 $T=210000 42560 0 0 $X=209570 $Y=41920
X8590 1 2 867 874 DLY1JI3VX1 $T=215600 51520 0 0 $X=215170 $Y=50880
X8591 1 2 1094 99 DLY1JI3VX1 $T=217840 42560 1 0 $X=217410 $Y=37440
X8592 1 2 1078 1325 DLY1JI3VX1 $T=217840 60480 1 0 $X=217410 $Y=55360
X8593 1 2 1253 1254 DLY1JI3VX1 $T=231840 33600 0 0 $X=231410 $Y=32960
X8594 1 2 443 1255 DLY1JI3VX1 $T=231840 42560 0 0 $X=231410 $Y=41920
X8595 1 2 1326 1092 DLY1JI3VX1 $T=234080 168000 1 0 $X=233650 $Y=162880
X8596 1 2 1260 1328 DLY1JI3VX1 $T=235200 168000 0 0 $X=234770 $Y=167360
X8597 1 2 1174 721 DLY1JI3VX1 $T=236320 150080 1 0 $X=235890 $Y=144960
X8598 1 2 863 450 DLY1JI3VX1 $T=238000 141120 1 0 $X=237570 $Y=136000
X8599 1 2 884 1259 DLY1JI3VX1 $T=244160 33600 0 0 $X=243730 $Y=32960
X8600 1 2 458 1104 DLY1JI3VX1 $T=245280 141120 1 0 $X=244850 $Y=136000
X8601 1 2 1097 1262 DLY1JI3VX1 $T=246960 33600 1 0 $X=246530 $Y=28480
X8602 1 2 1271 1108 DLY1JI3VX1 $T=253120 78400 0 0 $X=252690 $Y=77760
X8603 1 2 1106 1266 DLY1JI3VX1 $T=254240 42560 0 0 $X=253810 $Y=41920
X8604 1 2 482 1110 DLY1JI3VX1 $T=255360 159040 0 0 $X=254930 $Y=158400
X8605 1 2 491 1270 DLY1JI3VX1 $T=260960 42560 0 0 $X=260530 $Y=41920
X8606 1 2 722 1274 DLY1JI3VX1 $T=265440 150080 1 0 $X=265010 $Y=144960
X8607 1 2 502 1275 DLY1JI3VX1 $T=266560 42560 0 0 $X=266130 $Y=41920
X8608 1 2 1117 1119 DLY1JI3VX1 $T=270480 168000 1 0 $X=270050 $Y=162880
X8609 1 2 1264 1120 DLY1JI3VX1 $T=272160 132160 0 0 $X=271730 $Y=131520
X8610 1 2 723 1278 DLY1JI3VX1 $T=273840 42560 0 0 $X=273410 $Y=41920
X8611 1 2 1276 1279 DLY1JI3VX1 $T=277760 150080 0 0 $X=277330 $Y=149440
X8612 1 2 724 1121 DLY1JI3VX1 $T=283920 69440 0 0 $X=283490 $Y=68800
X8613 1 2 533 916 DLY1JI3VX1 $T=286160 168000 0 0 $X=285730 $Y=167360
X8614 1 2 530 101 DLY1JI3VX1 $T=288400 114240 0 0 $X=287970 $Y=113600
X8615 1 2 1122 1282 DLY1JI3VX1 $T=289520 42560 0 0 $X=289090 $Y=41920
X8616 1 2 915 1124 DLY1JI3VX1 $T=289520 69440 0 0 $X=289090 $Y=68800
X8617 1 2 918 1283 DLY1JI3VX1 $T=293440 159040 1 0 $X=293010 $Y=153920
X8618 1 2 1284 1285 DLY1JI3VX1 $T=297920 42560 0 0 $X=297490 $Y=41920
X8619 1 2 725 1287 DLY1JI3VX1 $T=303520 42560 0 0 $X=303090 $Y=41920
X8620 1 2 547 552 DLY1JI3VX1 $T=303520 159040 1 0 $X=303090 $Y=153920
X8621 1 2 551 1288 DLY1JI3VX1 $T=304640 33600 0 0 $X=304210 $Y=32960
X8622 1 2 726 1290 DLY1JI3VX1 $T=309120 42560 0 0 $X=308690 $Y=41920
X8623 1 2 1301 1291 DLY1JI3VX1 $T=309680 159040 0 0 $X=309250 $Y=158400
X8624 1 2 727 1292 DLY1JI3VX1 $T=315280 42560 0 0 $X=314850 $Y=41920
X8625 1 2 578 1337 DLY1JI3VX1 $T=316400 159040 1 0 $X=315970 $Y=153920
X8626 1 2 728 1294 DLY1JI3VX1 $T=320880 42560 0 0 $X=320450 $Y=41920
X8627 1 2 1129 595 DLY1JI3VX1 $T=327040 42560 1 0 $X=326610 $Y=37440
X8628 1 2 1296 596 DLY1JI3VX1 $T=327040 60480 0 0 $X=326610 $Y=59840
X8629 1 2 644 1299 DLY1JI3VX1 $T=336000 42560 1 180 $X=329970 $Y=41920
X8630 1 2 1137 1304 DLY1JI3VX1 $T=336000 42560 0 0 $X=335570 $Y=41920
X8631 1 2 940 1338 DLY1JI3VX1 $T=337680 141120 0 0 $X=337250 $Y=140480
X8632 1 2 979 1305 DLY1JI3VX1 $T=347760 176960 0 180 $X=341730 $Y=171840
X8633 1 2 729 625 DLY1JI3VX1 $T=342720 51520 0 0 $X=342290 $Y=50880
X8634 1 2 1136 1141 DLY1JI3VX1 $T=352240 60480 0 180 $X=346210 $Y=55360
X8635 1 2 980 620 DLY1JI3VX1 $T=352240 141120 1 180 $X=346210 $Y=140480
X8636 1 2 731 1147 DLY1JI3VX1 $T=360080 150080 1 0 $X=359650 $Y=144960
X8637 1 2 1310 1150 DLY1JI3VX1 $T=364560 168000 0 0 $X=364130 $Y=167360
X8638 1 2 733 1151 DLY1JI3VX1 $T=365680 150080 1 0 $X=365250 $Y=144960
X8639 1 2 1155 957 DLY1JI3VX1 $T=371840 33600 0 0 $X=371410 $Y=32960
X8640 1 2 942 1153 DLY1JI3VX1 $T=379120 141120 0 180 $X=373090 $Y=136000
X8641 1 2 956 651 DLY1JI3VX1 $T=373520 159040 0 0 $X=373090 $Y=158400
X8642 1 2 1154 1311 DLY1JI3VX1 $T=374080 33600 1 0 $X=373650 $Y=28480
X8643 1 2 941 654 DLY1JI3VX1 $T=374080 132160 0 0 $X=373650 $Y=131520
X8644 1 2 734 660 DLY1JI3VX1 $T=375200 185920 1 0 $X=374770 $Y=180800
X8645 1 2 1163 144 DLY1JI3VX1 $T=379680 33600 0 0 $X=379250 $Y=32960
X8646 1 2 964 1340 DLY1JI3VX1 $T=385840 24640 1 0 $X=385410 $Y=19520
X8647 1 2 963 1313 DLY1JI3VX1 $T=388640 33600 1 0 $X=388210 $Y=28480
X8648 1 2 686 1164 DLY1JI3VX1 $T=389760 78400 1 0 $X=389330 $Y=73280
X8649 1 2 698 699 DLY1JI3VX1 $T=407680 33600 0 0 $X=407250 $Y=32960
X8650 1 2 737 700 DLY1JI3VX1 $T=413280 42560 0 0 $X=412850 $Y=41920
X8651 1 2 975 701 DLY1JI3VX1 $T=413280 51520 1 0 $X=412850 $Y=46400
X8652 1 2 738 702 DLY1JI3VX1 $T=413280 51520 0 0 $X=412850 $Y=50880
X8653 1 2 222 422 374 397 415 OR4JI3VX1 $T=184240 24640 0 0 $X=183810 $Y=24000
X8654 1 2 484 451 386 460 353 OR4JI3VX1 $T=199920 24640 0 180 $X=193330 $Y=19520
X8655 1 2 409 405 858 499 419 OR4JI3VX1 $T=206080 24640 0 0 $X=205650 $Y=24000
X8656 1 2 1148 634 1316 953 944 OR4JI3VX1 $T=366800 24640 1 180 $X=360210 $Y=24000
X8657 1 2 154 739 84 150 DFRRQJI3VX1 $T=21280 176960 1 0 $X=20850 $Y=171840
X8658 1 2 154 147 84 160 DFRRQJI3VX1 $T=21840 159040 0 0 $X=21410 $Y=158400
X8659 1 2 154 148 84 157 DFRRQJI3VX1 $T=21840 185920 1 0 $X=21410 $Y=180800
X8660 1 2 154 982 84 153 DFRRQJI3VX1 $T=22400 150080 1 0 $X=21970 $Y=144960
X8661 1 2 154 149 84 162 DFRRQJI3VX1 $T=22960 194880 1 0 $X=22530 $Y=189760
X8662 1 2 154 155 84 146 DFRRQJI3VX1 $T=39200 105280 0 180 $X=23650 $Y=100160
X8663 1 2 154 164 84 703 DFRRQJI3VX1 $T=39760 105280 1 180 $X=24210 $Y=104640
X8664 1 2 154 191 84 704 DFRRQJI3VX1 $T=39760 114240 0 180 $X=24210 $Y=109120
X8665 1 2 154 741 84 745 DFRRQJI3VX1 $T=24640 123200 0 0 $X=24210 $Y=122560
X8666 1 2 154 740 84 747 DFRRQJI3VX1 $T=24640 132160 1 0 $X=24210 $Y=127040
X8667 1 2 154 984 84 746 DFRRQJI3VX1 $T=24640 132160 0 0 $X=24210 $Y=131520
X8668 1 2 154 990 84 756 DFRRQJI3VX1 $T=39200 150080 1 0 $X=38770 $Y=144960
X8669 1 2 154 193 84 158 DFRRQJI3VX1 $T=54880 114240 1 180 $X=39330 $Y=113600
X8670 1 2 154 743 84 751 DFRRQJI3VX1 $T=39760 141120 1 0 $X=39330 $Y=136000
X8671 1 2 154 744 84 752 DFRRQJI3VX1 $T=39760 141120 0 0 $X=39330 $Y=140480
X8672 1 2 154 171 84 173 DFRRQJI3VX1 $T=39760 194880 1 0 $X=39330 $Y=189760
X8673 1 2 154 181 84 159 DFRRQJI3VX1 $T=56000 123200 0 180 $X=40450 $Y=118080
X8674 1 2 154 177 84 987 DFRRQJI3VX1 $T=57120 132160 0 180 $X=41570 $Y=127040
X8675 1 2 154 1181 84 1182 DFRRQJI3VX1 $T=42000 132160 0 0 $X=41570 $Y=131520
X8676 1 2 180 1179 84 779 DFRRQJI3VX1 $T=44800 42560 1 0 $X=44370 $Y=37440
X8677 1 2 180 1183 84 762 DFRRQJI3VX1 $T=44800 42560 0 0 $X=44370 $Y=41920
X8678 1 2 180 166 84 187 DFRRQJI3VX1 $T=44800 51520 1 0 $X=44370 $Y=46400
X8679 1 2 180 190 84 705 DFRRQJI3VX1 $T=44800 51520 0 0 $X=44370 $Y=50880
X8680 1 2 180 748 84 709 DFRRQJI3VX1 $T=45360 60480 1 0 $X=44930 $Y=55360
X8681 1 2 180 749 84 185 DFRRQJI3VX1 $T=45920 69440 1 0 $X=45490 $Y=64320
X8682 1 2 154 1185 84 753 DFRRQJI3VX1 $T=62720 194880 1 180 $X=47170 $Y=194240
X8683 1 2 154 86 84 708 DFRRQJI3VX1 $T=50960 203840 1 0 $X=50530 $Y=198720
X8684 1 2 154 188 84 768 DFRRQJI3VX1 $T=57120 141120 1 0 $X=56690 $Y=136000
X8685 1 2 154 1194 84 759 DFRRQJI3VX1 $T=72240 141120 1 180 $X=56690 $Y=140480
X8686 1 2 154 1000 84 201 DFRRQJI3VX1 $T=72240 150080 0 180 $X=56690 $Y=144960
X8687 1 2 154 200 84 203 DFRRQJI3VX1 $T=58240 203840 0 0 $X=57810 $Y=203200
X8688 1 2 180 1192 84 773 DFRRQJI3VX1 $T=62160 51520 1 0 $X=61730 $Y=46400
X8689 1 2 180 189 84 1003 DFRRQJI3VX1 $T=62160 60480 1 0 $X=61730 $Y=55360
X8690 1 2 180 1187 84 223 DFRRQJI3VX1 $T=62720 42560 1 0 $X=62290 $Y=37440
X8691 1 2 180 1190 84 776 DFRRQJI3VX1 $T=62720 42560 0 0 $X=62290 $Y=41920
X8692 1 2 180 997 84 218 DFRRQJI3VX1 $T=63280 60480 0 0 $X=62850 $Y=59840
X8693 1 2 180 112 84 710 DFRRQJI3VX1 $T=63840 51520 0 0 $X=63410 $Y=50880
X8694 1 2 154 769 84 780 DFRRQJI3VX1 $T=72240 168000 1 0 $X=71810 $Y=162880
X8695 1 2 154 235 84 1394 DFRRQJI3VX1 $T=87360 168000 1 180 $X=71810 $Y=167360
X8696 1 2 154 976 84 1193 DFRRQJI3VX1 $T=89040 141120 0 180 $X=73490 $Y=136000
X8697 1 2 154 1168 84 182 DFRRQJI3VX1 $T=89040 150080 0 180 $X=73490 $Y=144960
X8698 1 2 154 1318 84 772 DFRRQJI3VX1 $T=89600 203840 1 180 $X=74050 $Y=203200
X8699 1 2 154 229 84 215 DFRRQJI3VX1 $T=90160 185920 0 180 $X=74610 $Y=180800
X8700 1 2 154 261 84 782 DFRRQJI3VX1 $T=75040 212800 1 0 $X=74610 $Y=207680
X8701 1 2 154 230 84 1198 DFRRQJI3VX1 $T=75600 176960 1 0 $X=75170 $Y=171840
X8702 1 2 154 234 84 213 DFRRQJI3VX1 $T=90720 176960 1 180 $X=75170 $Y=176320
X8703 1 2 154 1005 84 212 DFRRQJI3VX1 $T=90720 194880 1 180 $X=75170 $Y=194240
X8704 1 2 180 224 84 1001 DFRRQJI3VX1 $T=78400 60480 0 0 $X=77970 $Y=59840
X8705 1 2 180 1196 84 232 DFRRQJI3VX1 $T=78960 51520 1 0 $X=78530 $Y=46400
X8706 1 2 180 774 84 783 DFRRQJI3VX1 $T=78960 51520 0 0 $X=78530 $Y=50880
X8707 1 2 180 1002 84 236 DFRRQJI3VX1 $T=78960 60480 1 0 $X=78530 $Y=55360
X8708 1 2 180 216 84 711 DFRRQJI3VX1 $T=100240 78400 1 180 $X=84690 $Y=77760
X8709 1 2 180 1200 84 712 DFRRQJI3VX1 $T=100240 141120 1 180 $X=84690 $Y=140480
X8710 1 2 154 239 84 225 DFRRQJI3VX1 $T=100240 194880 0 180 $X=84690 $Y=189760
X8711 1 2 154 1197 84 289 DFRRQJI3VX1 $T=100240 212800 1 180 $X=84690 $Y=212160
X8712 1 2 243 797 84 241 DFRRQJI3VX1 $T=98560 42560 1 0 $X=98130 $Y=37440
X8713 1 2 243 1209 84 245 DFRRQJI3VX1 $T=98560 42560 0 0 $X=98130 $Y=41920
X8714 1 2 180 233 84 792 DFRRQJI3VX1 $T=98560 51520 1 0 $X=98130 $Y=46400
X8715 1 2 180 1008 84 242 DFRRQJI3VX1 $T=98560 51520 0 0 $X=98130 $Y=50880
X8716 1 2 180 1007 84 1009 DFRRQJI3VX1 $T=98560 60480 1 0 $X=98130 $Y=55360
X8717 1 2 180 770 84 1199 DFRRQJI3VX1 $T=98560 60480 0 0 $X=98130 $Y=59840
X8718 1 2 154 217 84 789 DFRRQJI3VX1 $T=98560 150080 1 0 $X=98130 $Y=144960
X8719 1 2 154 237 84 788 DFRRQJI3VX1 $T=98560 168000 0 0 $X=98130 $Y=167360
X8720 1 2 244 240 84 246 DFRRQJI3VX1 $T=98560 194880 0 0 $X=98130 $Y=194240
X8721 1 2 247 1201 84 821 DFRRQJI3VX1 $T=98560 212800 1 0 $X=98130 $Y=207680
X8722 1 2 248 1214 84 117 DFRRQJI3VX1 $T=100240 212800 0 0 $X=99810 $Y=212160
X8723 1 2 180 262 84 1202 DFRRQJI3VX1 $T=102480 123200 1 0 $X=102050 $Y=118080
X8724 1 2 180 1205 84 256 DFRRQJI3VX1 $T=103040 132160 0 0 $X=102610 $Y=131520
X8725 1 2 255 1010 98 1011 DFRRQJI3VX1 $T=103600 150080 0 0 $X=103170 $Y=149440
X8726 1 2 257 771 84 1204 DFRRQJI3VX1 $T=104160 176960 1 0 $X=103730 $Y=171840
X8727 1 2 258 1012 84 808 DFRRQJI3VX1 $T=104720 141120 1 0 $X=104290 $Y=136000
X8728 1 2 154 795 84 260 DFRRQJI3VX1 $T=104720 176960 0 0 $X=104290 $Y=176320
X8729 1 2 1013 271 84 798 DFRRQJI3VX1 $T=108640 203840 0 0 $X=108210 $Y=203200
X8730 1 2 154 781 84 264 DFRRQJI3VX1 $T=109760 194880 1 0 $X=109330 $Y=189760
X8731 1 2 243 785 84 252 DFRRQJI3VX1 $T=128800 51520 1 180 $X=113250 $Y=50880
X8732 1 2 243 276 84 791 DFRRQJI3VX1 $T=128800 60480 0 180 $X=113250 $Y=55360
X8733 1 2 243 249 84 800 DFRRQJI3VX1 $T=113680 60480 0 0 $X=113250 $Y=59840
X8734 1 2 154 714 84 1016 DFRRQJI3VX1 $T=113680 194880 0 0 $X=113250 $Y=194240
X8735 1 2 243 1031 84 268 DFRRQJI3VX1 $T=114240 42560 1 0 $X=113810 $Y=37440
X8736 1 2 243 277 84 802 DFRRQJI3VX1 $T=114240 42560 0 0 $X=113810 $Y=41920
X8737 1 2 243 1206 84 790 DFRRQJI3VX1 $T=129360 51520 0 180 $X=113810 $Y=46400
X8738 1 2 243 1022 84 801 DFRRQJI3VX1 $T=114800 33600 0 0 $X=114370 $Y=32960
X8739 1 2 180 259 84 1360 DFRRQJI3VX1 $T=118160 114240 0 0 $X=117730 $Y=113600
X8740 1 2 180 799 84 1203 DFRRQJI3VX1 $T=133280 123200 0 180 $X=117730 $Y=118080
X8741 1 2 180 275 84 715 DFRRQJI3VX1 $T=119840 132160 0 0 $X=119410 $Y=131520
X8742 1 2 180 265 84 296 DFRRQJI3VX1 $T=119840 141120 1 0 $X=119410 $Y=136000
X8743 1 2 180 266 98 1017 DFRRQJI3VX1 $T=119840 150080 0 0 $X=119410 $Y=149440
X8744 1 2 280 1023 84 806 DFRRQJI3VX1 $T=119840 176960 0 0 $X=119410 $Y=176320
X8745 1 2 285 270 84 1018 DFRRQJI3VX1 $T=121520 176960 1 0 $X=121090 $Y=171840
X8746 1 2 287 1208 84 1019 DFRRQJI3VX1 $T=122080 168000 0 0 $X=121650 $Y=167360
X8747 1 2 180 1027 84 329 DFRRQJI3VX1 $T=123200 132160 1 0 $X=122770 $Y=127040
X8748 1 2 243 293 92 273 DFRRQJI3VX1 $T=145600 105280 0 180 $X=130050 $Y=100160
X8749 1 2 243 811 92 299 DFRRQJI3VX1 $T=131040 51520 1 0 $X=130610 $Y=46400
X8750 1 2 243 1039 92 279 DFRRQJI3VX1 $T=146160 51520 1 180 $X=130610 $Y=50880
X8751 1 2 243 1041 92 288 DFRRQJI3VX1 $T=146160 60480 0 180 $X=130610 $Y=55360
X8752 1 2 243 283 92 1034 DFRRQJI3VX1 $T=131040 60480 0 0 $X=130610 $Y=59840
X8753 1 2 243 1021 92 1032 DFRRQJI3VX1 $T=131040 69440 1 0 $X=130610 $Y=64320
X8754 1 2 243 1220 92 817 DFRRQJI3VX1 $T=131600 42560 0 0 $X=131170 $Y=41920
X8755 1 2 180 807 92 284 DFRRQJI3VX1 $T=148960 114240 0 180 $X=133410 $Y=109120
X8756 1 2 180 1215 98 307 DFRRQJI3VX1 $T=134960 141120 0 0 $X=134530 $Y=140480
X8757 1 2 180 294 98 302 DFRRQJI3VX1 $T=135520 159040 1 0 $X=135090 $Y=153920
X8758 1 2 180 88 98 337 DFRRQJI3VX1 $T=136080 141120 1 0 $X=135650 $Y=136000
X8759 1 2 255 1211 98 291 DFRRQJI3VX1 $T=136080 176960 0 0 $X=135650 $Y=176320
X8760 1 2 255 1212 98 1030 DFRRQJI3VX1 $T=136640 194880 1 0 $X=136210 $Y=189760
X8761 1 2 306 89 98 1217 DFRRQJI3VX1 $T=138320 203840 0 0 $X=137890 $Y=203200
X8762 1 2 243 327 92 1026 DFRRQJI3VX1 $T=160160 96320 1 180 $X=144610 $Y=95680
X8763 1 2 243 1319 92 1045 DFRRQJI3VX1 $T=145600 69440 0 0 $X=145170 $Y=68800
X8764 1 2 243 1042 92 1033 DFRRQJI3VX1 $T=160720 105280 0 180 $X=145170 $Y=100160
X8765 1 2 243 311 92 1048 DFRRQJI3VX1 $T=147280 69440 1 0 $X=146850 $Y=64320
X8766 1 2 243 1222 92 322 DFRRQJI3VX1 $T=147840 42560 0 0 $X=147410 $Y=41920
X8767 1 2 243 1226 92 1036 DFRRQJI3VX1 $T=162960 51520 0 180 $X=147410 $Y=46400
X8768 1 2 243 1049 92 813 DFRRQJI3VX1 $T=162960 51520 1 180 $X=147410 $Y=50880
X8769 1 2 243 1225 92 812 DFRRQJI3VX1 $T=162960 60480 1 180 $X=147410 $Y=59840
X8770 1 2 180 822 98 321 DFRRQJI3VX1 $T=151200 159040 1 0 $X=150770 $Y=153920
X8771 1 2 180 1223 98 820 DFRRQJI3VX1 $T=166320 168000 1 180 $X=150770 $Y=167360
X8772 1 2 255 815 98 118 DFRRQJI3VX1 $T=166320 176960 1 180 $X=150770 $Y=176320
X8773 1 2 180 1224 98 309 DFRRQJI3VX1 $T=166880 150080 0 180 $X=151330 $Y=144960
X8774 1 2 306 336 98 1058 DFRRQJI3VX1 $T=151760 185920 1 0 $X=151330 $Y=180800
X8775 1 2 306 338 98 1053 DFRRQJI3VX1 $T=152320 185920 0 0 $X=151890 $Y=185280
X8776 1 2 306 339 98 364 DFRRQJI3VX1 $T=152320 194880 1 0 $X=151890 $Y=189760
X8777 1 2 306 1050 98 316 DFRRQJI3VX1 $T=170800 203840 1 180 $X=155250 $Y=203200
X8778 1 2 243 1054 92 825 DFRRQJI3VX1 $T=173600 105280 1 180 $X=158050 $Y=104640
X8779 1 2 243 1046 98 335 DFRRQJI3VX1 $T=159040 132160 0 0 $X=158610 $Y=131520
X8780 1 2 243 831 92 1004 DFRRQJI3VX1 $T=175840 105280 0 180 $X=160290 $Y=100160
X8781 1 2 306 331 98 355 DFRRQJI3VX1 $T=160720 212800 0 0 $X=160290 $Y=212160
X8782 1 2 243 829 92 1052 DFRRQJI3VX1 $T=176960 96320 1 180 $X=161410 $Y=95680
X8783 1 2 243 326 92 1059 DFRRQJI3VX1 $T=163520 69440 1 0 $X=163090 $Y=64320
X8784 1 2 243 1227 92 323 DFRRQJI3VX1 $T=179200 42560 0 180 $X=163650 $Y=37440
X8785 1 2 243 1233 92 342 DFRRQJI3VX1 $T=179760 42560 1 180 $X=164210 $Y=41920
X8786 1 2 243 325 92 836 DFRRQJI3VX1 $T=164640 60480 1 0 $X=164210 $Y=55360
X8787 1 2 243 1229 92 334 DFRRQJI3VX1 $T=180320 51520 0 180 $X=164770 $Y=46400
X8788 1 2 243 841 92 1228 DFRRQJI3VX1 $T=165200 51520 0 0 $X=164770 $Y=50880
X8789 1 2 180 93 98 333 DFRRQJI3VX1 $T=181440 168000 0 180 $X=165890 $Y=162880
X8790 1 2 180 1057 98 350 DFRRQJI3VX1 $T=183120 159040 0 180 $X=167570 $Y=153920
X8791 1 2 243 1231 92 819 DFRRQJI3VX1 $T=188160 114240 0 180 $X=172610 $Y=109120
X8792 1 2 243 1064 98 349 DFRRQJI3VX1 $T=189840 132160 1 180 $X=174290 $Y=131520
X8793 1 2 243 1239 92 828 DFRRQJI3VX1 $T=190400 105280 1 180 $X=174850 $Y=104640
X8794 1 2 243 843 92 356 DFRRQJI3VX1 $T=190960 105280 0 180 $X=175410 $Y=100160
X8795 1 2 306 1063 98 379 DFRRQJI3VX1 $T=176960 212800 0 0 $X=176530 $Y=212160
X8796 1 2 243 1323 98 847 DFRRQJI3VX1 $T=193200 141120 1 180 $X=177650 $Y=140480
X8797 1 2 243 1237 92 365 DFRRQJI3VX1 $T=197120 42560 1 180 $X=181570 $Y=41920
X8798 1 2 243 1240 92 121 DFRRQJI3VX1 $T=197680 51520 0 180 $X=182130 $Y=46400
X8799 1 2 243 366 92 383 DFRRQJI3VX1 $T=182560 51520 0 0 $X=182130 $Y=50880
X8800 1 2 243 838 92 1072 DFRRQJI3VX1 $T=182560 60480 1 0 $X=182130 $Y=55360
X8801 1 2 243 403 92 348 DFRRQJI3VX1 $T=197680 123200 0 180 $X=182130 $Y=118080
X8802 1 2 387 1235 98 368 DFRRQJI3VX1 $T=197680 150080 0 180 $X=182130 $Y=144960
X8803 1 2 387 1241 98 361 DFRRQJI3VX1 $T=198240 150080 1 180 $X=182690 $Y=149440
X8804 1 2 243 1242 92 367 DFRRQJI3VX1 $T=198800 114240 1 180 $X=183250 $Y=113600
X8805 1 2 387 1345 98 407 DFRRQJI3VX1 $T=183680 159040 1 0 $X=183250 $Y=153920
X8806 1 2 387 1362 98 839 DFRRQJI3VX1 $T=184240 168000 1 0 $X=183810 $Y=162880
X8807 1 2 243 875 92 717 DFRRQJI3VX1 $T=203280 87360 1 180 $X=187730 $Y=86720
X8808 1 2 243 392 92 375 DFRRQJI3VX1 $T=203280 96320 0 180 $X=187730 $Y=91200
X8809 1 2 243 396 92 1066 DFRRQJI3VX1 $T=203280 114240 0 180 $X=187730 $Y=109120
X8810 1 2 243 1075 98 373 DFRRQJI3VX1 $T=203280 123200 1 180 $X=187730 $Y=122560
X8811 1 2 243 95 98 1234 DFRRQJI3VX1 $T=203280 132160 0 180 $X=187730 $Y=127040
X8812 1 2 406 1324 98 859 DFRRQJI3VX1 $T=192640 168000 0 0 $X=192210 $Y=167360
X8813 1 2 306 1245 98 395 DFRRQJI3VX1 $T=208320 212800 0 180 $X=192770 $Y=207680
X8814 1 2 387 388 98 1326 DFRRQJI3VX1 $T=198240 150080 1 0 $X=197810 $Y=144960
X8815 1 2 387 389 98 1174 DFRRQJI3VX1 $T=198240 150080 0 0 $X=197810 $Y=149440
X8816 1 2 387 1074 92 867 DFRRQJI3VX1 $T=199920 69440 1 0 $X=199490 $Y=64320
X8817 1 2 243 404 92 394 DFRRQJI3VX1 $T=215040 114240 1 180 $X=199490 $Y=113600
X8818 1 2 243 424 92 398 DFRRQJI3VX1 $T=215600 51520 0 180 $X=200050 $Y=46400
X8819 1 2 243 874 92 402 DFRRQJI3VX1 $T=215600 51520 1 180 $X=200050 $Y=50880
X8820 1 2 387 377 92 719 DFRRQJI3VX1 $T=201040 60480 0 0 $X=200610 $Y=59840
X8821 1 2 441 1325 92 413 DFRRQJI3VX1 $T=202720 60480 1 0 $X=202290 $Y=55360
X8822 1 2 871 1363 98 97 DFRRQJI3VX1 $T=204400 176960 0 0 $X=203970 $Y=176320
X8823 1 2 387 371 92 1078 DFRRQJI3VX1 $T=223440 69440 1 180 $X=207890 $Y=68800
X8824 1 2 306 1089 98 1080 DFRRQJI3VX1 $T=225680 212800 0 180 $X=210130 $Y=207680
X8825 1 2 387 860 98 863 DFRRQJI3VX1 $T=228480 141120 0 180 $X=212930 $Y=136000
X8826 1 2 387 1249 98 1082 DFRRQJI3VX1 $T=228480 141120 1 180 $X=212930 $Y=140480
X8827 1 2 387 1115 98 1056 DFRRQJI3VX1 $T=228480 150080 0 180 $X=212930 $Y=144960
X8828 1 2 868 455 98 1083 DFRRQJI3VX1 $T=228480 150080 1 180 $X=212930 $Y=149440
X8829 1 2 441 1328 98 1071 DFRRQJI3VX1 $T=228480 159040 1 180 $X=212930 $Y=158400
X8830 1 2 441 99 92 862 DFRRQJI3VX1 $T=226800 42560 1 0 $X=226370 $Y=37440
X8831 1 2 441 1254 92 444 DFRRQJI3VX1 $T=226800 51520 1 0 $X=226370 $Y=46400
X8832 1 2 441 1255 92 428 DFRRQJI3VX1 $T=226800 51520 0 0 $X=226370 $Y=50880
X8833 1 2 441 877 92 443 DFRRQJI3VX1 $T=226800 60480 1 0 $X=226370 $Y=55360
X8834 1 2 441 1087 92 1253 DFRRQJI3VX1 $T=226800 60480 0 0 $X=226370 $Y=59840
X8835 1 2 441 430 92 1094 DFRRQJI3VX1 $T=226800 69440 1 0 $X=226370 $Y=64320
X8836 1 2 442 1251 98 133 DFRRQJI3VX1 $T=226800 176960 0 0 $X=226370 $Y=176320
X8837 1 2 442 1329 98 888 DFRRQJI3VX1 $T=226800 185920 1 0 $X=226370 $Y=180800
X8838 1 2 442 1252 98 1095 DFRRQJI3VX1 $T=226800 194880 1 0 $X=226370 $Y=189760
X8839 1 2 442 876 98 1090 DFRRQJI3VX1 $T=226800 203840 0 0 $X=226370 $Y=203200
X8840 1 2 442 436 98 440 DFRRQJI3VX1 $T=229600 212800 1 0 $X=229170 $Y=207680
X8841 1 2 442 1092 98 886 DFRRQJI3VX1 $T=230720 159040 1 0 $X=230290 $Y=153920
X8842 1 2 442 721 98 446 DFRRQJI3VX1 $T=231280 150080 0 0 $X=230850 $Y=149440
X8843 1 2 442 450 98 1103 DFRRQJI3VX1 $T=232960 141120 0 0 $X=232530 $Y=140480
X8844 1 2 457 438 92 458 DFRRQJI3VX1 $T=236320 114240 1 0 $X=235890 $Y=109120
X8845 1 2 454 872 98 722 DFRRQJI3VX1 $T=236880 132160 0 0 $X=236450 $Y=131520
X8846 1 2 441 1259 92 461 DFRRQJI3VX1 $T=239120 42560 0 0 $X=238690 $Y=41920
X8847 1 2 457 445 98 1264 DFRRQJI3VX1 $T=240240 123200 0 0 $X=239810 $Y=122560
X8848 1 2 457 1104 98 895 DFRRQJI3VX1 $T=240240 132160 1 0 $X=239810 $Y=127040
X8849 1 2 442 1332 98 892 DFRRQJI3VX1 $T=240240 203840 1 0 $X=239810 $Y=198720
X8850 1 2 441 1262 92 471 DFRRQJI3VX1 $T=241920 42560 1 0 $X=241490 $Y=37440
X8851 1 2 441 1266 92 1096 DFRRQJI3VX1 $T=257040 51520 0 180 $X=241490 $Y=46400
X8852 1 2 441 878 92 1106 DFRRQJI3VX1 $T=241920 51520 0 0 $X=241490 $Y=50880
X8853 1 2 441 1108 92 881 DFRRQJI3VX1 $T=257040 60480 0 180 $X=241490 $Y=55360
X8854 1 2 441 434 92 1097 DFRRQJI3VX1 $T=257040 60480 1 180 $X=241490 $Y=59840
X8855 1 2 441 879 92 884 DFRRQJI3VX1 $T=257040 69440 0 180 $X=241490 $Y=64320
X8856 1 2 442 1333 98 456 DFRRQJI3VX1 $T=259840 203840 1 180 $X=244290 $Y=203200
X8857 1 2 442 1274 98 459 DFRRQJI3VX1 $T=261520 150080 1 180 $X=245970 $Y=149440
X8858 1 2 442 1110 98 453 DFRRQJI3VX1 $T=261520 159040 0 180 $X=245970 $Y=153920
X8859 1 2 442 1265 98 479 DFRRQJI3VX1 $T=249200 212800 1 0 $X=248770 $Y=207680
X8860 1 2 442 465 98 1260 DFRRQJI3VX1 $T=265440 150080 0 180 $X=249890 $Y=144960
X8861 1 2 441 1107 92 1271 DFRRQJI3VX1 $T=252000 69440 0 0 $X=251570 $Y=68800
X8862 1 2 457 1120 98 476 DFRRQJI3VX1 $T=272160 132160 0 180 $X=256610 $Y=127040
X8863 1 2 441 1275 92 475 DFRRQJI3VX1 $T=272720 51520 0 180 $X=257170 $Y=46400
X8864 1 2 441 1278 92 497 DFRRQJI3VX1 $T=257600 51520 0 0 $X=257170 $Y=50880
X8865 1 2 441 509 92 502 DFRRQJI3VX1 $T=257600 60480 0 0 $X=257170 $Y=59840
X8866 1 2 441 896 92 723 DFRRQJI3VX1 $T=272720 69440 0 180 $X=257170 $Y=64320
X8867 1 2 441 1270 92 501 DFRRQJI3VX1 $T=258160 60480 1 0 $X=257730 $Y=55360
X8868 1 2 457 510 98 1276 DFRRQJI3VX1 $T=259280 123200 0 0 $X=258850 $Y=122560
X8869 1 2 457 449 92 1117 DFRRQJI3VX1 $T=259840 123200 1 0 $X=259410 $Y=118080
X8870 1 2 442 1119 98 493 DFRRQJI3VX1 $T=276080 159040 1 180 $X=260530 $Y=158400
X8871 1 2 442 1273 98 490 DFRRQJI3VX1 $T=276080 203840 1 180 $X=260530 $Y=203200
X8872 1 2 442 1279 98 1268 DFRRQJI3VX1 $T=277200 159040 0 180 $X=261650 $Y=153920
X8873 1 2 442 503 98 482 DFRRQJI3VX1 $T=277760 150080 1 180 $X=262210 $Y=149440
X8874 1 2 441 489 92 491 DFRRQJI3VX1 $T=282240 69440 1 180 $X=266690 $Y=68800
X8875 1 2 441 1121 92 512 DFRRQJI3VX1 $T=291200 51520 0 180 $X=275650 $Y=46400
X8876 1 2 441 1282 92 517 DFRRQJI3VX1 $T=291200 51520 1 180 $X=275650 $Y=50880
X8877 1 2 441 1124 92 516 DFRRQJI3VX1 $T=291200 60480 0 180 $X=275650 $Y=55360
X8878 1 2 441 504 92 1122 DFRRQJI3VX1 $T=276080 60480 0 0 $X=275650 $Y=59840
X8879 1 2 441 1277 92 915 DFRRQJI3VX1 $T=276080 69440 1 0 $X=275650 $Y=64320
X8880 1 2 441 513 92 724 DFRRQJI3VX1 $T=276640 96320 1 0 $X=276210 $Y=91200
X8881 1 2 457 101 98 127 DFRRQJI3VX1 $T=291760 123200 0 180 $X=276210 $Y=118080
X8882 1 2 457 911 98 530 DFRRQJI3VX1 $T=277200 123200 0 0 $X=276770 $Y=122560
X8883 1 2 442 908 98 100 DFRRQJI3VX1 $T=292320 194880 1 180 $X=276770 $Y=194240
X8884 1 2 457 538 98 918 DFRRQJI3VX1 $T=277760 159040 0 0 $X=277330 $Y=158400
X8885 1 2 457 520 98 533 DFRRQJI3VX1 $T=278320 159040 1 0 $X=277890 $Y=153920
X8886 1 2 442 1283 98 518 DFRRQJI3VX1 $T=293440 168000 0 180 $X=277890 $Y=162880
X8887 1 2 442 916 98 909 DFRRQJI3VX1 $T=295120 176960 0 180 $X=279570 $Y=171840
X8888 1 2 442 912 98 506 DFRRQJI3VX1 $T=295120 194880 0 180 $X=279570 $Y=189760
X8889 1 2 457 565 102 547 DFRRQJI3VX1 $T=292320 150080 0 0 $X=291890 $Y=149440
X8890 1 2 441 1285 92 532 DFRRQJI3VX1 $T=309120 51520 0 180 $X=293570 $Y=46400
X8891 1 2 441 1290 92 920 DFRRQJI3VX1 $T=309120 51520 1 180 $X=293570 $Y=50880
X8892 1 2 441 1287 92 531 DFRRQJI3VX1 $T=309120 60480 0 180 $X=293570 $Y=55360
X8893 1 2 441 1127 92 1284 DFRRQJI3VX1 $T=294000 60480 0 0 $X=293570 $Y=59840
X8894 1 2 441 558 92 725 DFRRQJI3VX1 $T=294000 69440 1 0 $X=293570 $Y=64320
X8895 1 2 457 552 102 426 DFRRQJI3VX1 $T=309120 159040 1 180 $X=293570 $Y=158400
X8896 1 2 441 562 92 726 DFRRQJI3VX1 $T=294560 78400 1 0 $X=294130 $Y=73280
X8897 1 2 441 1288 92 1125 DFRRQJI3VX1 $T=310240 42560 0 180 $X=294690 $Y=37440
X8898 1 2 441 563 92 551 DFRRQJI3VX1 $T=295120 69440 0 0 $X=294690 $Y=68800
X8899 1 2 590 923 116 555 DFRRQJI3VX1 $T=297360 212800 1 0 $X=296930 $Y=207680
X8900 1 2 457 921 102 578 DFRRQJI3VX1 $T=307440 150080 0 0 $X=307010 $Y=149440
X8901 1 2 441 1294 102 560 DFRRQJI3VX1 $T=326480 51520 0 180 $X=310930 $Y=46400
X8902 1 2 441 1292 102 137 DFRRQJI3VX1 $T=326480 51520 1 180 $X=310930 $Y=50880
X8903 1 2 441 596 102 570 DFRRQJI3VX1 $T=326480 60480 0 180 $X=310930 $Y=55360
X8904 1 2 441 607 102 1129 DFRRQJI3VX1 $T=326480 69440 0 180 $X=310930 $Y=64320
X8905 1 2 457 1336 102 591 DFRRQJI3VX1 $T=311360 185920 1 0 $X=310930 $Y=180800
X8906 1 2 441 595 102 1134 DFRRQJI3VX1 $T=311920 42560 1 0 $X=311490 $Y=37440
X8907 1 2 441 606 102 728 DFRRQJI3VX1 $T=327040 60480 1 180 $X=311490 $Y=59840
X8908 1 2 441 602 102 1296 DFRRQJI3VX1 $T=311920 69440 0 0 $X=311490 $Y=68800
X8909 1 2 441 571 102 727 DFRRQJI3VX1 $T=311920 78400 1 0 $X=311490 $Y=73280
X8910 1 2 457 1128 102 589 DFRRQJI3VX1 $T=311920 185920 0 0 $X=311490 $Y=185280
X8911 1 2 590 1131 116 559 DFRRQJI3VX1 $T=327600 203840 1 180 $X=312050 $Y=203200
X8912 1 2 590 569 116 576 DFRRQJI3VX1 $T=314720 203840 1 0 $X=314290 $Y=198720
X8913 1 2 457 1295 102 940 DFRRQJI3VX1 $T=322000 132160 1 0 $X=321570 $Y=127040
X8914 1 2 457 572 102 941 DFRRQJI3VX1 $T=322000 132160 0 0 $X=321570 $Y=131520
X8915 1 2 457 930 102 1301 DFRRQJI3VX1 $T=322000 141120 1 0 $X=321570 $Y=136000
X8916 1 2 457 1338 102 585 DFRRQJI3VX1 $T=337120 150080 0 180 $X=321570 $Y=144960
X8917 1 2 457 1337 102 609 DFRRQJI3VX1 $T=322000 159040 1 0 $X=321570 $Y=153920
X8918 1 2 457 573 102 733 DFRRQJI3VX1 $T=322560 141120 0 0 $X=322130 $Y=140480
X8919 1 2 457 574 102 942 DFRRQJI3VX1 $T=322560 150080 0 0 $X=322130 $Y=149440
X8920 1 2 457 1291 102 580 DFRRQJI3VX1 $T=338240 159040 1 180 $X=322690 $Y=158400
X8921 1 2 441 1304 102 592 DFRRQJI3VX1 $T=342720 51520 0 180 $X=327170 $Y=46400
X8922 1 2 441 625 102 594 DFRRQJI3VX1 $T=342720 51520 1 180 $X=327170 $Y=50880
X8923 1 2 441 629 102 1137 DFRRQJI3VX1 $T=328160 60480 1 0 $X=327730 $Y=55360
X8924 1 2 441 628 102 729 DFRRQJI3VX1 $T=328160 69440 1 0 $X=327730 $Y=64320
X8925 1 2 457 604 102 600 DFRRQJI3VX1 $T=329280 185920 0 0 $X=328850 $Y=185280
X8926 1 2 457 1300 102 139 DFRRQJI3VX1 $T=329840 194880 0 0 $X=329410 $Y=194240
X8927 1 2 590 1353 116 730 DFRRQJI3VX1 $T=336000 203840 0 0 $X=335570 $Y=203200
X8928 1 2 457 103 102 979 DFRRQJI3VX1 $T=355040 132160 0 180 $X=339490 $Y=127040
X8929 1 2 457 1305 102 608 DFRRQJI3VX1 $T=355040 150080 1 180 $X=339490 $Y=149440
X8930 1 2 457 620 102 617 DFRRQJI3VX1 $T=355040 159040 0 180 $X=339490 $Y=153920
X8931 1 2 457 597 102 731 DFRRQJI3VX1 $T=355600 132160 1 180 $X=340050 $Y=131520
X8932 1 2 457 1153 102 674 DFRRQJI3VX1 $T=355600 141120 0 180 $X=340050 $Y=136000
X8933 1 2 457 1147 102 610 DFRRQJI3VX1 $T=355600 150080 0 180 $X=340050 $Y=144960
X8934 1 2 457 1299 102 616 DFRRQJI3VX1 $T=356720 42560 1 180 $X=341170 $Y=41920
X8935 1 2 457 635 102 1136 DFRRQJI3VX1 $T=356720 60480 1 180 $X=341170 $Y=59840
X8936 1 2 457 1141 102 1149 DFRRQJI3VX1 $T=355040 51520 0 0 $X=354610 $Y=50880
X8937 1 2 105 952 102 644 DFRRQJI3VX1 $T=355040 69440 1 0 $X=354610 $Y=64320
X8938 1 2 105 631 102 636 DFRRQJI3VX1 $T=355040 194880 1 0 $X=354610 $Y=189760
X8939 1 2 105 1306 102 630 DFRRQJI3VX1 $T=355040 194880 0 0 $X=354610 $Y=194240
X8940 1 2 105 656 102 956 DFRRQJI3VX1 $T=357280 150080 0 0 $X=356850 $Y=149440
X8941 1 2 105 657 102 980 DFRRQJI3VX1 $T=357840 159040 1 0 $X=357410 $Y=153920
X8942 1 2 105 1308 102 1310 DFRRQJI3VX1 $T=358400 141120 1 0 $X=357970 $Y=136000
X8943 1 2 105 1151 102 662 DFRRQJI3VX1 $T=358400 141120 0 0 $X=357970 $Y=140480
X8944 1 2 105 651 102 950 DFRRQJI3VX1 $T=358400 159040 0 0 $X=357970 $Y=158400
X8945 1 2 105 1150 102 1142 DFRRQJI3VX1 $T=358400 168000 1 0 $X=357970 $Y=162880
X8946 1 2 105 654 102 659 DFRRQJI3VX1 $T=358960 132160 0 0 $X=358530 $Y=131520
X8947 1 2 457 1311 102 732 DFRRQJI3VX1 $T=377440 42560 1 180 $X=361890 $Y=41920
X8948 1 2 105 1157 102 1154 DFRRQJI3VX1 $T=362320 60480 0 0 $X=361890 $Y=59840
X8949 1 2 457 957 102 143 DFRRQJI3VX1 $T=378000 51520 0 180 $X=362450 $Y=46400
X8950 1 2 105 655 102 1155 DFRRQJI3VX1 $T=362880 60480 1 0 $X=362450 $Y=55360
X8951 1 2 105 660 102 642 DFRRQJI3VX1 $T=380800 176960 1 180 $X=365250 $Y=176320
X8952 1 2 105 1158 102 734 DFRRQJI3VX1 $T=381360 176960 0 180 $X=365810 $Y=171840
X8953 1 2 105 959 102 646 DFRRQJI3VX1 $T=388640 150080 1 180 $X=373090 $Y=149440
X8954 1 2 105 144 102 650 DFRRQJI3VX1 $T=394800 51520 0 180 $X=379250 $Y=46400
X8955 1 2 105 1340 102 647 DFRRQJI3VX1 $T=395360 42560 0 180 $X=379810 $Y=37440
X8956 1 2 105 1313 102 653 DFRRQJI3VX1 $T=395360 42560 1 180 $X=379810 $Y=41920
X8957 1 2 105 1164 102 645 DFRRQJI3VX1 $T=395360 51520 1 180 $X=379810 $Y=50880
X8958 1 2 105 736 102 963 DFRRQJI3VX1 $T=380240 60480 1 0 $X=379810 $Y=55360
X8959 1 2 105 735 102 686 DFRRQJI3VX1 $T=380240 60480 0 0 $X=379810 $Y=59840
X8960 1 2 105 958 102 964 DFRRQJI3VX1 $T=380240 69440 1 0 $X=379810 $Y=64320
X8961 1 2 105 666 102 1163 DFRRQJI3VX1 $T=380240 69440 0 0 $X=379810 $Y=68800
X8962 1 2 105 970 102 683 DFRRQJI3VX1 $T=408800 150080 1 180 $X=393250 $Y=149440
X8963 1 2 105 965 102 681 DFRRQJI3VX1 $T=409920 132160 0 180 $X=394370 $Y=127040
X8964 1 2 105 699 102 694 DFRRQJI3VX1 $T=413280 42560 0 180 $X=397730 $Y=37440
X8965 1 2 105 700 102 971 DFRRQJI3VX1 $T=413280 42560 1 180 $X=397730 $Y=41920
X8966 1 2 105 701 102 691 DFRRQJI3VX1 $T=413280 51520 0 180 $X=397730 $Y=46400
X8967 1 2 105 702 102 689 DFRRQJI3VX1 $T=413280 51520 1 180 $X=397730 $Y=50880
X8968 1 2 105 692 102 738 DFRRQJI3VX1 $T=398160 60480 1 0 $X=397730 $Y=55360
X8969 1 2 105 1167 102 737 DFRRQJI3VX1 $T=398160 60480 0 0 $X=397730 $Y=59840
X8970 1 2 105 106 102 975 DFRRQJI3VX1 $T=398160 69440 1 0 $X=397730 $Y=64320
X8971 1 2 105 107 102 698 DFRRQJI3VX1 $T=398160 69440 0 0 $X=397730 $Y=68800
X8972 1 2 105 108 102 521 DFRRQJI3VX1 $T=398160 105280 1 0 $X=397730 $Y=100160
X8973 1 2 153 167 INJI3VX1 $T=42000 159040 1 0 $X=41570 $Y=153920
X8974 1 2 162 988 INJI3VX1 $T=42560 176960 0 0 $X=42130 $Y=176320
X8975 1 2 173 991 INJI3VX1 $T=50960 176960 0 0 $X=50530 $Y=176320
X8976 1 2 708 192 INJI3VX1 $T=63840 194880 1 0 $X=63410 $Y=189760
X8977 1 2 231 1062 INJI3VX1 $T=181440 150080 0 0 $X=181010 $Y=149440
X8978 1 2 127 220 INJI3VX1 $T=202720 176960 0 0 $X=202290 $Y=176320
X8979 1 2 231 1091 INJI3VX1 $T=231840 176960 1 0 $X=231410 $Y=171840
X8980 1 2 1091 442 INJI3VX1 $T=233520 168000 0 0 $X=233090 $Y=167360
X8981 1 2 440 1093 INJI3VX1 $T=238560 203840 1 0 $X=238130 $Y=198720
X8982 1 2 892 893 INJI3VX1 $T=247520 185920 0 0 $X=247090 $Y=185280
X8983 1 2 123 590 INJI3VX1 $T=309120 203840 0 0 $X=308690 $Y=203200
X8984 1 2 681 668 INJI3VX1 $T=392560 132160 1 0 $X=392130 $Y=127040
X8985 1 2 1062 180 INJI3VX2 $T=180320 150080 1 0 $X=179890 $Y=144960
X8986 1 2 206 DAC<1> BUJI3VX12 $T=69440 24640 0 180 $X=56690 $Y=19520
X8987 1 2 777 DAC<2> BUJI3VX12 $T=77840 24640 1 180 $X=65090 $Y=24000
X8988 1 2 778 DAC<3> BUJI3VX12 $T=82880 24640 0 180 $X=70130 $Y=19520
X8989 1 2 160 163 147 983 151 ON22JI3VX1 $T=33600 159040 0 180 $X=28690 $Y=153920
X8990 1 2 157 985 1395 156 150 ON22JI3VX1 $T=36400 168000 1 180 $X=31490 $Y=167360
X8991 1 2 745 161 750 988 747 ON22JI3VX1 $T=40320 168000 1 0 $X=39890 $Y=162880
X8992 1 2 707 1390 1185 178 1184 ON22JI3VX1 $T=58800 185920 1 180 $X=53890 $Y=185280
X8993 1 2 759 192 1189 1188 1394 ON22JI3VX1 $T=63280 168000 0 0 $X=62850 $Y=167360
X8994 1 2 1188 219 200 178 205 ON22JI3VX1 $T=71680 194880 0 180 $X=66770 $Y=189760
X8995 1 2 1331 485 1329 1100 448 ON22JI3VX1 $T=246400 185920 0 180 $X=241490 $Y=180800
X8996 1 2 462 485 1333 1263 472 ON22JI3VX1 $T=251440 194880 1 0 $X=251010 $Y=189760
X8997 1 2 493 492 898 1112 1268 ON22JI3VX1 $T=267680 185920 1 180 $X=262770 $Y=185280
X8998 1 2 585 931 564 1132 580 ON22JI3VX1 $T=319760 159040 1 180 $X=314850 $Y=158400
X8999 1 2 600 612 1302 946 139 ON22JI3VX1 $T=344960 185920 0 180 $X=340050 $Y=180800
X9000 1 2 642 1146 603 104 1142 ON22JI3VX1 $T=364560 168000 1 180 $X=359650 $Y=167360
X9001 1 2 690 687 676 672 693 ON22JI3VX1 $T=392560 114240 0 180 $X=387650 $Y=109120
X9002 1 2 695 966 970 981 683 ON22JI3VX1 $T=398720 159040 1 0 $X=398290 $Y=153920
X9003 1 2 1236 391 851 124 400 AN31JI3VX1 $T=195440 185920 0 0 $X=195010 $Y=185280
X9004 1 2 487 1113 894 1272 505 AN31JI3VX1 $T=264320 168000 0 0 $X=263890 $Y=167360
X9005 1 2 1396 1289 1351 549 1286 AN31JI3VX1 $T=313040 168000 0 180 $X=308690 $Y=162880
X9006 1 2 1359 202 1397 1189 NO3JI3VX0 $T=63840 176960 1 0 $X=63410 $Y=171840
X9007 1 2 1380 1376 1098 452 NO3JI3VX0 $T=246400 159040 0 0 $X=245970 $Y=158400
X9008 1 2 534 542 1398 550 NO3JI3VX0 $T=295120 212800 0 0 $X=294690 $Y=212160
X9009 1 2 220 587 136 925 NO3JI3VX0 $T=305200 176960 0 0 $X=304770 $Y=176320
X9010 1 2 381 386 196 858 410 OR4JI3VX2 $T=194320 24640 0 0 $X=193890 $Y=24000
X9011 1 2 1169 289 117 282 HAJI3VX1 $T=138320 203840 1 180 $X=130050 $Y=203200
X9012 1 2 1399 289 316 816 HAJI3VX1 $T=158480 212800 0 180 $X=150210 $Y=207680
X9013 1 2 834 343 1058 347 HAJI3VX1 $T=175840 185920 0 180 $X=167570 $Y=180800
X9014 1 2 352 1055 355 835 HAJI3VX1 $T=173600 203840 0 0 $X=173170 $Y=203200
X9015 1 2 1400 1053 347 362 HAJI3VX1 $T=175280 185920 0 0 $X=174850 $Y=185280
X9016 1 2 845 379 835 128 HAJI3VX1 $T=186480 203840 0 0 $X=186050 $Y=203200
X9017 1 2 480 479 1401 474 HAJI3VX1 $T=262080 194880 1 180 $X=253810 $Y=194240
X9018 1 2 486 490 474 483 HAJI3VX1 $T=267680 203840 0 180 $X=259410 $Y=198720
X9019 1 2 569 576 932 566 HAJI3VX1 $T=316960 212800 1 0 $X=316530 $Y=207680
X9020 1 2 583 1123 589 1297 HAJI3VX1 $T=322000 176960 0 0 $X=321570 $Y=176320
X9021 1 2 1135 593 1402 932 HAJI3VX1 $T=329840 212800 0 0 $X=329410 $Y=212160
X9022 1 2 1143 630 945 1145 HAJI3VX1 $T=351680 176960 1 180 $X=343410 $Y=176320
X9023 1 2 1269 437 DLY4JI3VX1 $T=252000 212800 0 0 $X=251570 $Y=212160
X9024 1 2 755 1374 176 NO2I1JI3VX1 $T=50400 150080 0 0 $X=49970 $Y=149440
X9025 1 2 819 303 302 NO2I1JI3VX1 $T=143360 123200 0 0 $X=142930 $Y=122560
X9026 1 2 828 320 321 NO2I1JI3VX1 $T=166320 132160 0 180 $X=162530 $Y=127040
X9027 1 2 368 122 1053 NO2I1JI3VX1 $T=184240 185920 0 0 $X=183810 $Y=185280
X9028 1 2 1053 1070 368 NO2I1JI3VX1 $T=187600 185920 0 0 $X=187170 $Y=185280
X9029 1 2 376 94 378 NO2I1JI3VX1 $T=187600 203840 1 0 $X=187170 $Y=198720
X9030 1 2 407 390 426 NO2I1JI3VX1 $T=197680 176960 1 0 $X=197250 $Y=171840
X9031 1 2 857 304 129 NO2I1JI3VX1 $T=202720 168000 0 180 $X=198930 $Y=162880
X9032 1 2 855 418 414 NO2I1JI3VX1 $T=210000 159040 0 180 $X=206210 $Y=153920
X9033 1 2 1090 96 426 NO2I1JI3VX1 $T=219520 194880 1 180 $X=215730 $Y=194240
X9034 1 2 426 1088 1090 NO2I1JI3VX1 $T=235200 194880 1 180 $X=231410 $Y=194240
X9035 1 2 889 464 466 NO2I1JI3VX1 $T=249760 168000 1 0 $X=249330 $Y=162880
X9036 1 2 909 505 506 NO2I1JI3VX1 $T=278320 176960 0 180 $X=274530 $Y=171840
X9037 1 2 515 905 518 NO2I1JI3VX1 $T=280560 168000 1 180 $X=276770 $Y=167360
X9038 1 2 542 1130 553 NO2I1JI3VX1 $T=306880 123200 0 0 $X=306450 $Y=122560
X9039 1 2 582 1352 580 NO2I1JI3VX1 $T=332640 168000 0 180 $X=328850 $Y=162880
X9040 1 2 608 599 600 NO2I1JI3VX1 $T=337120 176960 0 180 $X=333330 $Y=171840
X9041 1 2 600 928 608 NO2I1JI3VX1 $T=338800 168000 1 180 $X=335010 $Y=167360
X9042 1 2 152 1395 169 150 739 AO22JI3VX1 $T=31360 168000 1 180 $X=25890 $Y=167360
X9043 1 2 170 152 162 220 149 AO22JI3VX1 $T=44240 185920 1 180 $X=38770 $Y=185280
X9044 1 2 754 152 993 220 171 AO22JI3VX1 $T=50960 185920 1 180 $X=45490 $Y=185280
X9045 1 2 773 318 227 223 221 AO22JI3VX1 $T=86800 42560 0 180 $X=81330 $Y=37440
X9046 1 2 236 318 227 779 222 AO22JI3VX1 $T=89040 33600 0 180 $X=83570 $Y=28480
X9047 1 2 776 318 227 762 429 AO22JI3VX1 $T=95200 33600 0 180 $X=89730 $Y=28480
X9048 1 2 232 318 227 783 451 AO22JI3VX1 $T=103040 33600 0 0 $X=102610 $Y=32960
X9049 1 2 242 318 227 241 484 AO22JI3VX1 $T=109760 33600 0 0 $X=109330 $Y=32960
X9050 1 2 252 318 227 245 405 AO22JI3VX1 $T=112000 33600 1 0 $X=111570 $Y=28480
X9051 1 2 1024 313 310 798 271 AO22JI3VX1 $T=130480 203840 1 180 $X=125010 $Y=203200
X9052 1 2 268 318 227 801 409 AO22JI3VX1 $T=126560 24640 0 0 $X=126130 $Y=24000
X9053 1 2 803 313 310 296 265 AO22JI3VX1 $T=131600 141120 1 180 $X=126130 $Y=140480
X9054 1 2 804 313 310 1017 266 AO22JI3VX1 $T=132160 159040 0 180 $X=126690 $Y=153920
X9055 1 2 1014 313 310 1018 270 AO22JI3VX1 $T=132160 185920 0 180 $X=126690 $Y=180800
X9056 1 2 1028 313 310 1016 714 AO22JI3VX1 $T=133840 194880 1 180 $X=128370 $Y=194240
X9057 1 2 272 313 310 1019 1208 AO22JI3VX1 $T=129360 168000 1 0 $X=128930 $Y=162880
X9058 1 2 1169 313 310 117 1214 AO22JI3VX1 $T=137760 212800 1 0 $X=137330 $Y=207680
X9059 1 2 814 319 125 291 1211 AO22JI3VX1 $T=146160 168000 1 180 $X=140690 $Y=167360
X9060 1 2 292 319 125 118 815 AO22JI3VX1 $T=141680 185920 1 0 $X=141250 $Y=180800
X9061 1 2 1040 319 125 1030 1212 AO22JI3VX1 $T=146720 194880 1 180 $X=141250 $Y=194240
X9062 1 2 279 318 227 288 415 AO22JI3VX1 $T=142240 33600 0 0 $X=141810 $Y=32960
X9063 1 2 1029 319 125 1217 89 AO22JI3VX1 $T=143360 212800 1 0 $X=142930 $Y=207680
X9064 1 2 1219 319 125 302 294 AO22JI3VX1 $T=150640 159040 1 180 $X=145170 $Y=158400
X9065 1 2 299 318 227 817 422 AO22JI3VX1 $T=148960 24640 0 0 $X=148530 $Y=24000
X9066 1 2 308 319 125 321 822 AO22JI3VX1 $T=150640 159040 0 0 $X=150210 $Y=158400
X9067 1 2 313 827 310 309 1224 AO22JI3VX1 $T=155120 141120 1 0 $X=154690 $Y=136000
X9068 1 2 812 318 227 1036 397 AO22JI3VX1 $T=156240 33600 0 0 $X=155810 $Y=32960
X9069 1 2 319 330 125 820 1223 AO22JI3VX1 $T=163520 159040 1 180 $X=158050 $Y=158400
X9070 1 2 313 1320 310 335 1046 AO22JI3VX1 $T=165760 141120 0 180 $X=160290 $Y=136000
X9071 1 2 1399 319 125 340 1050 AO22JI3VX1 $T=160720 212800 1 0 $X=160290 $Y=207680
X9072 1 2 323 318 227 322 460 AO22JI3VX1 $T=163520 33600 1 0 $X=163090 $Y=28480
X9073 1 2 319 830 125 333 93 AO22JI3VX1 $T=166880 159040 0 0 $X=166450 $Y=158400
X9074 1 2 834 313 310 1058 336 AO22JI3VX1 $T=174160 176960 1 180 $X=168690 $Y=176320
X9075 1 2 1400 313 310 1053 338 AO22JI3VX1 $T=174160 185920 1 180 $X=168690 $Y=185280
X9076 1 2 1403 313 310 364 339 AO22JI3VX1 $T=174160 194880 0 180 $X=168690 $Y=189760
X9077 1 2 352 319 125 355 331 AO22JI3VX1 $T=174160 212800 0 180 $X=168690 $Y=207680
X9078 1 2 342 318 227 334 353 AO22JI3VX1 $T=170240 24640 0 0 $X=169810 $Y=24000
X9079 1 2 319 1343 125 350 1057 AO22JI3VX1 $T=181440 159040 1 180 $X=175970 $Y=158400
X9080 1 2 313 837 310 349 1064 AO22JI3VX1 $T=180320 141120 1 0 $X=179890 $Y=136000
X9081 1 2 845 319 125 379 1063 AO22JI3VX1 $T=187040 212800 0 180 $X=181570 $Y=207680
X9082 1 2 365 318 227 121 499 AO22JI3VX1 $T=187040 33600 0 0 $X=186610 $Y=32960
X9083 1 2 1404 319 125 395 1245 AO22JI3VX1 $T=201040 203840 0 0 $X=200610 $Y=203200
X9084 1 2 402 318 227 398 419 AO22JI3VX1 $T=205520 42560 1 0 $X=205090 $Y=37440
X9085 1 2 480 1170 1256 479 1265 AO22JI3VX1 $T=260960 194880 0 180 $X=255490 $Y=189760
X9086 1 2 478 473 898 902 1114 AO22JI3VX1 $T=259840 176960 0 0 $X=259410 $Y=176320
X9087 1 2 486 1170 1256 490 1273 AO22JI3VX1 $T=262640 194880 0 0 $X=262210 $Y=194240
X9088 1 2 475 488 447 497 634 AO22JI3VX1 $T=266560 33600 1 0 $X=266130 $Y=28480
X9089 1 2 507 1170 1256 100 908 AO22JI3VX1 $T=270480 194880 0 0 $X=270050 $Y=194240
X9090 1 2 531 488 447 532 924 AO22JI3VX1 $T=299040 33600 1 0 $X=298610 $Y=28480
X9091 1 2 583 587 925 589 1128 AO22JI3VX1 $T=314720 194880 0 180 $X=309250 $Y=189760
X9092 1 2 579 587 925 591 1336 AO22JI3VX1 $T=320880 176960 1 180 $X=315410 $Y=176320
X9093 1 2 570 488 447 137 632 AO22JI3VX1 $T=320320 33600 0 0 $X=319890 $Y=32960
X9094 1 2 560 488 447 1134 934 AO22JI3VX1 $T=320880 33600 1 0 $X=320450 $Y=28480
X9095 1 2 139 598 587 1302 1300 AO22JI3VX1 $T=341600 194880 0 180 $X=336130 $Y=189760
X9096 1 2 1143 587 925 630 1306 AO22JI3VX1 $T=352240 185920 1 180 $X=346770 $Y=185280
X9097 1 2 196 pulse_active BUJI3VX6 $T=55440 24640 0 0 $X=55010 $Y=24000
X9098 1 2 775 116 BUJI3VX6 $T=77280 123200 0 0 $X=76850 $Y=122560
X9099 1 2 1405 457 BUJI3VX6 $T=285600 132160 0 0 $X=285170 $Y=131520
X9100 1 2 646 447 BUJI3VX6 $T=373520 150080 1 0 $X=373090 $Y=144960
X9101 1 2 153 151 163 982 1406 ON31JI3VX1 $T=32480 150080 1 180 $X=27570 $Y=149440
X9102 1 2 157 986 178 148 1407 ON31JI3VX1 $T=36960 176960 1 180 $X=32050 $Y=176320
X9103 1 2 708 199 178 86 763 ON31JI3VX1 $T=63840 194880 0 180 $X=58930 $Y=189760
X9104 1 2 839 360 358 1362 1344 ON31JI3VX1 $T=180320 168000 0 0 $X=179890 $Y=167360
X9105 1 2 1080 416 1347 1089 1248 ON31JI3VX1 $T=211120 203840 0 0 $X=210690 $Y=203200
X9106 1 2 892 1258 485 1332 1257 ON31JI3VX1 $T=249760 194880 1 180 $X=244850 $Y=194240
X9107 1 2 506 903 485 912 910 ON31JI3VX1 $T=274400 194880 1 0 $X=273970 $Y=189760
X9108 1 2 1297 1293 1352 581 586 ON31JI3VX1 $T=328720 168000 1 180 $X=323810 $Y=167360
X9109 1 2 600 601 948 604 938 ON31JI3VX1 $T=331520 185920 1 0 $X=331090 $Y=180800
X9110 1 2 636 947 948 631 641 ON31JI3VX1 $T=347200 194880 1 0 $X=346770 $Y=189760
X9111 1 2 681 1312 145 965 1408 ON31JI3VX1 $T=392000 123200 1 0 $X=391570 $Y=118080
X9112 1 2 1159 966 981 969 967 ON31JI3VX1 $T=394800 168000 1 0 $X=394370 $Y=162880
X9113 1 2 337 349 354 837 EO3JI3VX1 $T=167440 141120 0 0 $X=167010 $Y=140480
X9114 1 2 337 350 359 1343 EO3JI3VX1 $T=169680 150080 1 0 $X=169250 $Y=144960
X9115 1 2 231 154 BUJI3VX2 $T=124880 194880 1 0 $X=124450 $Y=189760
X9116 1 2 380 417 BUJI3VX2 $T=192640 212800 0 0 $X=192210 $Y=212160
X9117 1 2 447 227 BUJI3VX2 $T=216160 33600 0 0 $X=215730 $Y=32960
X9118 1 2 431 231 BUJI3VX2 $T=220640 185920 1 0 $X=220210 $Y=180800
X9119 1 2 488 318 BUJI3VX2 $T=241920 33600 1 180 $X=238130 $Y=32960
X9120 1 2 494 267 BUJI3VX2 $T=268800 212800 1 180 $X=265010 $Y=212160
X9121 1 2 525 1405 BUJI3VX2 $T=282240 132160 0 0 $X=281810 $Y=131520
X9122 1 2 540 554 BUJI3VX2 $T=305760 203840 0 0 $X=305330 $Y=203200
X9123 1 2 588 up_switches<16> BUJI3VX2 $T=328160 24640 1 0 $X=327730 $Y=19520
X9124 1 2 584 up_switches<17> BUJI3VX2 $T=332080 24640 1 0 $X=331650 $Y=19520
X9125 1 2 605 up_switches<18> BUJI3VX2 $T=335440 24640 1 0 $X=335010 $Y=19520
X9126 1 2 917 up_switches<19> BUJI3VX2 $T=342720 24640 1 0 $X=342290 $Y=19520
X9127 1 2 924 up_switches<21> BUJI3VX2 $T=352240 24640 1 180 $X=348450 $Y=24000
X9128 1 2 634 up_switches<20> BUJI3VX2 $T=362880 24640 0 180 $X=359090 $Y=19520
X9129 1 2 632 up_switches<23> BUJI3VX2 $T=360640 33600 1 0 $X=360210 $Y=28480
X9130 1 2 953 up_switches<26> BUJI3VX2 $T=362880 24640 1 0 $X=362450 $Y=19520
X9131 1 2 944 up_switches<25> BUJI3VX2 $T=366800 24640 0 0 $X=366370 $Y=24000
X9132 1 2 934 up_switches<24> BUJI3VX2 $T=366800 33600 1 0 $X=366370 $Y=28480
X9133 1 2 1148 up_switches<27> BUJI3VX2 $T=370160 24640 0 0 $X=369730 $Y=24000
X9134 1 2 457 105 BUJI3VX2 $T=372960 51520 0 0 $X=372530 $Y=50880
X9135 1 2 658 up_switches<28> BUJI3VX2 $T=381360 24640 1 0 $X=380930 $Y=19520
X9136 1 2 652 up_switches<29> BUJI3VX2 $T=397600 24640 0 180 $X=393810 $Y=19520
X9137 1 2 1160 up_switches<30> BUJI3VX2 $T=402640 24640 0 180 $X=398850 $Y=19520
X9138 1 2 697 up_switches<31> BUJI3VX2 $T=402640 24640 1 0 $X=402210 $Y=19520
X9139 1 2 220 enable INJI3VX3 $T=92960 176960 0 0 $X=92530 $Y=176320
X9140 1 2 1062 243 INJI3VX3 $T=181440 159040 0 0 $X=181010 $Y=158400
X9141 1 2 318 716 INJI3VX3 $T=194880 33600 1 0 $X=194450 $Y=28480
X9142 1 2 1409 900 INJI3VX3 $T=215600 212800 0 0 $X=215170 $Y=212160
X9143 1 2 1091 441 INJI3VX3 $T=233520 159040 1 180 $X=230290 $Y=158400
X9144 1 2 545 up_switches<14> INJI3VX3 $T=303520 24640 1 0 $X=303090 $Y=19520
X9145 1 2 548 up_switches<15> INJI3VX3 $T=308560 24640 1 0 $X=308130 $Y=19520
X9146 1 2 978 up_switches<22> INJI3VX3 $T=325920 24640 0 0 $X=325490 $Y=24000
X9147 1 2 869 220 1116 1246 NA3I2JI3VX1 $T=216160 168000 1 180 $X=211810 $Y=167360
X9148 1 2 96 1088 873 1346 NA3I2JI3VX1 $T=220640 194880 0 180 $X=216290 $Y=189760
X9149 1 2 556 559 555 550 NA3I2JI3VX1 $T=311920 212800 1 180 $X=307570 $Y=212160
X9150 1 2 603 599 586 1410 NA3I2JI3VX1 $T=334880 168000 1 180 $X=330530 $Y=167360
X9151 1 2 373 350 1051 832 EN3JI3VX1 $T=183120 123200 1 180 $X=172050 $Y=122560
X9152 1 2 115 748 154 183 109 748 SDFRRQJI3VX1 $T=62160 78400 1 180 $X=41570 $Y=77760
X9153 1 2 111 166 154 209 109 166 SDFRRQJI3VX1 $T=62160 96320 0 180 $X=41570 $Y=91200
X9154 1 2 113 155 154 253 109 155 SDFRRQJI3VX1 $T=62160 96320 1 180 $X=41570 $Y=95680
X9155 1 2 115 189 154 207 109 189 SDFRRQJI3VX1 $T=62720 69440 1 180 $X=42130 $Y=68800
X9156 1 2 111 190 154 207 109 190 SDFRRQJI3VX1 $T=62720 78400 0 180 $X=42130 $Y=73280
X9157 1 2 111 749 154 183 109 749 SDFRRQJI3VX1 $T=62720 87360 0 180 $X=42130 $Y=82240
X9158 1 2 113 164 154 204 109 164 SDFRRQJI3VX1 $T=62720 105280 0 180 $X=42130 $Y=100160
X9159 1 2 113 191 154 184 109 191 SDFRRQJI3VX1 $T=62720 105280 1 180 $X=42130 $Y=104640
X9160 1 2 113 193 154 251 109 193 SDFRRQJI3VX1 $T=63280 114240 0 180 $X=42690 $Y=109120
X9161 1 2 113 177 154 208 109 177 SDFRRQJI3VX1 $T=77280 123200 1 180 $X=56690 $Y=122560
X9162 1 2 113 181 154 254 109 181 SDFRRQJI3VX1 $T=80080 123200 0 180 $X=59490 $Y=118080
X9163 1 2 113 188 154 207 109 188 SDFRRQJI3VX1 $T=80080 132160 0 180 $X=59490 $Y=127040
X9164 1 2 115 112 180 208 109 112 SDFRRQJI3VX1 $T=64960 78400 0 0 $X=64530 $Y=77760
X9165 1 2 111 997 154 208 109 997 SDFRRQJI3VX1 $T=64960 87360 1 0 $X=64530 $Y=82240
X9166 1 2 115 224 154 209 109 224 SDFRRQJI3VX1 $T=64960 87360 0 0 $X=64530 $Y=86720
X9167 1 2 109 184 154 204 116 184 SDFRRQJI3VX1 $T=65520 96320 1 0 $X=65090 $Y=91200
X9168 1 2 109 204 154 208 116 204 SDFRRQJI3VX1 $T=65520 96320 0 0 $X=65090 $Y=95680
X9169 1 2 109 208 154 207 116 208 SDFRRQJI3VX1 $T=65520 105280 0 0 $X=65090 $Y=104640
X9170 1 2 109 207 154 183 116 207 SDFRRQJI3VX1 $T=66080 105280 1 0 $X=65650 $Y=100160
X9171 1 2 109 183 154 209 116 183 SDFRRQJI3VX1 $T=67760 114240 0 0 $X=67330 $Y=113600
X9172 1 2 113 230 154 209 109 230 SDFRRQJI3VX1 $T=70560 159040 1 0 $X=70130 $Y=153920
X9173 1 2 113 769 154 183 109 769 SDFRRQJI3VX1 $T=71120 150080 0 0 $X=70690 $Y=149440
X9174 1 2 111 233 180 204 109 233 SDFRRQJI3VX1 $T=95200 69440 0 180 $X=74610 $Y=64320
X9175 1 2 115 770 180 204 109 770 SDFRRQJI3VX1 $T=95200 69440 1 180 $X=74610 $Y=68800
X9176 1 2 115 216 180 184 109 216 SDFRRQJI3VX1 $T=95200 78400 0 180 $X=74610 $Y=73280
X9177 1 2 713 208 154 217 109 217 SDFRRQJI3VX1 $T=95200 114240 0 180 $X=74610 $Y=109120
X9178 1 2 113 976 154 250 109 976 SDFRRQJI3VX1 $T=95200 132160 1 180 $X=74610 $Y=131520
X9179 1 2 713 207 154 771 109 771 SDFRRQJI3VX1 $T=95200 159040 1 180 $X=74610 $Y=158400
X9180 1 2 109 253 154 184 116 253 SDFRRQJI3VX1 $T=103040 69440 1 0 $X=102610 $Y=64320
X9181 1 2 111 1007 180 184 109 1007 SDFRRQJI3VX1 $T=103040 78400 1 0 $X=102610 $Y=73280
X9182 1 2 713 204 180 262 109 262 SDFRRQJI3VX1 $T=103040 105280 1 0 $X=102610 $Y=100160
X9183 1 2 109 209 154 238 116 209 SDFRRQJI3VX1 $T=103040 123200 0 0 $X=102610 $Y=122560
X9184 1 2 713 184 180 1205 109 1205 SDFRRQJI3VX1 $T=103040 132160 1 0 $X=102610 $Y=127040
X9185 1 2 113 1200 180 332 109 1200 SDFRRQJI3VX1 $T=103040 141120 0 0 $X=102610 $Y=140480
X9186 1 2 113 237 154 238 109 237 SDFRRQJI3VX1 $T=103040 159040 1 0 $X=102610 $Y=153920
X9187 1 2 713 183 468 239 SPI_CS 239 SDFRRQJI3VX1 $T=103040 185920 1 0 $X=102610 $Y=180800
X9188 1 2 713 209 154 240 SPI_CS 240 SDFRRQJI3VX1 $T=103040 185920 0 0 $X=102610 $Y=185280
X9189 1 2 713 253 180 275 109 275 SDFRRQJI3VX1 $T=110320 105280 0 0 $X=109890 $Y=104640
X9190 1 2 115 276 243 253 109 276 SDFRRQJI3VX1 $T=110880 69440 0 0 $X=110450 $Y=68800
X9191 1 2 115 249 243 251 109 249 SDFRRQJI3VX1 $T=110880 87360 1 0 $X=110450 $Y=82240
X9192 1 2 111 277 243 251 109 277 SDFRRQJI3VX1 $T=110880 87360 0 0 $X=110450 $Y=86720
X9193 1 2 109 250 243 254 116 250 SDFRRQJI3VX1 $T=110880 96320 1 0 $X=110450 $Y=91200
X9194 1 2 111 1206 180 253 109 1206 SDFRRQJI3VX1 $T=111440 78400 0 0 $X=111010 $Y=77760
X9195 1 2 713 254 180 259 109 259 SDFRRQJI3VX1 $T=113680 114240 1 0 $X=113250 $Y=109120
X9196 1 2 713 238 468 261 SPI_CS 261 SDFRRQJI3VX1 $T=115360 212800 0 0 $X=114930 $Y=212160
X9197 1 2 109 251 180 253 116 251 SDFRRQJI3VX1 $T=123200 96320 0 0 $X=122770 $Y=95680
X9198 1 2 713 251 180 799 109 799 SDFRRQJI3VX1 $T=123200 123200 0 0 $X=122770 $Y=122560
X9199 1 2 111 1021 243 254 109 1021 SDFRRQJI3VX1 $T=131600 78400 1 0 $X=131170 $Y=73280
X9200 1 2 115 283 243 254 109 283 SDFRRQJI3VX1 $T=131600 87360 1 0 $X=131170 $Y=82240
X9201 1 2 109 254 180 251 116 254 SDFRRQJI3VX1 $T=132160 105280 0 0 $X=131730 $Y=104640
X9202 1 2 115 1319 243 238 109 1319 SDFRRQJI3VX1 $T=142240 96320 1 0 $X=141810 $Y=91200
X9203 1 2 111 1049 243 250 109 1049 SDFRRQJI3VX1 $T=142800 78400 0 0 $X=142370 $Y=77760
X9204 1 2 111 311 243 238 109 311 SDFRRQJI3VX1 $T=142800 87360 0 0 $X=142370 $Y=86720
X9205 1 2 343 310 231 313 98 343 SDFRRQJI3VX1 $T=149520 176960 1 0 $X=149090 $Y=171840
X9206 1 2 1055 125 231 319 98 1055 SDFRRQJI3VX1 $T=152880 194880 0 0 $X=152450 $Y=194240
X9207 1 2 115 325 243 332 109 325 SDFRRQJI3VX1 $T=162400 78400 1 0 $X=161970 $Y=73280
X9208 1 2 115 326 243 250 109 326 SDFRRQJI3VX1 $T=162400 87360 1 0 $X=161970 $Y=82240
X9209 1 2 111 841 243 332 109 841 SDFRRQJI3VX1 $T=162960 69440 0 0 $X=162530 $Y=68800
X9210 1 2 109 332 243 250 116 332 SDFRRQJI3VX1 $T=165760 87360 0 0 $X=165330 $Y=86720
X9211 1 2 113 829 243 370 109 829 SDFRRQJI3VX1 $T=186480 96320 0 180 $X=165890 $Y=91200
X9212 1 2 115 838 243 370 109 838 SDFRRQJI3VX1 $T=178640 60480 0 0 $X=178210 $Y=59840
X9213 1 2 111 366 243 370 109 366 SDFRRQJI3VX1 $T=179760 69440 1 0 $X=179330 $Y=64320
X9214 1 2 115 1074 468 372 109 1074 SDFRRQJI3VX1 $T=183120 78400 1 0 $X=182690 $Y=73280
X9215 1 2 111 371 468 854 109 371 SDFRRQJI3VX1 $T=203280 78400 1 180 $X=182690 $Y=77760
X9216 1 2 109 372 231 370 116 372 SDFRRQJI3VX1 $T=183120 96320 0 0 $X=182690 $Y=95680
X9217 1 2 109 370 231 332 116 370 SDFRRQJI3VX1 $T=187040 87360 1 0 $X=186610 $Y=82240
X9218 1 2 111 377 468 372 123 377 SDFRRQJI3VX1 $T=188160 69440 0 0 $X=187730 $Y=68800
X9219 1 2 713 370 468 860 SPI_CS 860 SDFRRQJI3VX1 $T=212240 141120 0 180 $X=191650 $Y=136000
X9220 1 2 713 250 468 388 SPI_CS 388 SDFRRQJI3VX1 $T=193200 141120 0 0 $X=192770 $Y=140480
X9221 1 2 713 332 468 389 SPI_CS 389 SDFRRQJI3VX1 $T=193200 159040 0 0 $X=192770 $Y=158400
X9222 1 2 115 1087 468 427 123 1087 SDFRRQJI3VX1 $T=223440 78400 0 180 $X=202850 $Y=73280
X9223 1 2 115 430 468 854 123 430 SDFRRQJI3VX1 $T=223440 78400 1 180 $X=202850 $Y=77760
X9224 1 2 113 875 468 854 123 875 SDFRRQJI3VX1 $T=223440 87360 1 180 $X=202850 $Y=86720
X9225 1 2 123 427 231 854 116 427 SDFRRQJI3VX1 $T=223440 96320 0 180 $X=202850 $Y=91200
X9226 1 2 123 854 231 372 116 854 SDFRRQJI3VX1 $T=223440 96320 1 180 $X=202850 $Y=95680
X9227 1 2 113 392 468 372 123 392 SDFRRQJI3VX1 $T=223440 105280 0 180 $X=202850 $Y=100160
X9228 1 2 113 396 468 427 123 396 SDFRRQJI3VX1 $T=223440 105280 1 180 $X=202850 $Y=104640
X9229 1 2 113 404 468 439 123 404 SDFRRQJI3VX1 $T=223440 114240 0 180 $X=202850 $Y=109120
X9230 1 2 113 95 468 435 123 95 SDFRRQJI3VX1 $T=223440 123200 1 180 $X=202850 $Y=122560
X9231 1 2 713 372 468 872 123 872 SDFRRQJI3VX1 $T=223440 132160 0 180 $X=202850 $Y=127040
X9232 1 2 113 1249 468 527 123 1249 SDFRRQJI3VX1 $T=223440 132160 1 180 $X=202850 $Y=131520
X9233 1 2 111 877 441 427 123 877 SDFRRQJI3VX1 $T=231840 69440 0 0 $X=231410 $Y=68800
X9234 1 2 123 238 442 437 116 238 SDFRRQJI3VX1 $T=231840 212800 0 0 $X=231410 $Y=212160
X9235 1 2 115 878 441 435 123 878 SDFRRQJI3VX1 $T=232960 78400 0 0 $X=232530 $Y=77760
X9236 1 2 111 434 441 439 123 434 SDFRRQJI3VX1 $T=232960 87360 1 0 $X=232530 $Y=82240
X9237 1 2 111 879 441 435 123 879 SDFRRQJI3VX1 $T=232960 87360 0 0 $X=232530 $Y=86720
X9238 1 2 123 439 441 427 116 439 SDFRRQJI3VX1 $T=232960 96320 0 0 $X=232530 $Y=95680
X9239 1 2 713 854 457 438 123 438 SDFRRQJI3VX1 $T=232960 105280 0 0 $X=232530 $Y=104640
X9240 1 2 123 435 457 439 116 435 SDFRRQJI3VX1 $T=233520 105280 1 0 $X=233090 $Y=100160
X9241 1 2 713 427 457 445 123 445 SDFRRQJI3VX1 $T=237440 114240 0 0 $X=237010 $Y=113600
X9242 1 2 713 435 457 449 123 449 SDFRRQJI3VX1 $T=239680 123200 1 0 $X=239250 $Y=118080
X9243 1 2 111 489 441 477 123 489 SDFRRQJI3VX1 $T=267680 78400 0 180 $X=247090 $Y=73280
X9244 1 2 113 1115 468 477 SPI_CS 1115 SDFRRQJI3VX1 $T=271040 141120 0 180 $X=250450 $Y=136000
X9245 1 2 113 455 442 514 SPI_CS 455 SDFRRQJI3VX1 $T=271040 141120 1 180 $X=250450 $Y=140480
X9246 1 2 113 465 457 526 SPI_CS 465 SDFRRQJI3VX1 $T=272160 132160 1 180 $X=251570 $Y=131520
X9247 1 2 115 1107 441 439 123 1107 SDFRRQJI3VX1 $T=254800 87360 1 0 $X=254370 $Y=82240
X9248 1 2 111 896 441 527 123 896 SDFRRQJI3VX1 $T=254800 87360 0 0 $X=254370 $Y=86720
X9249 1 2 115 509 441 527 123 509 SDFRRQJI3VX1 $T=255360 96320 1 0 $X=254930 $Y=91200
X9250 1 2 713 439 457 510 123 510 SDFRRQJI3VX1 $T=255920 114240 1 0 $X=255490 $Y=109120
X9251 1 2 123 477 441 435 116 477 SDFRRQJI3VX1 $T=256480 105280 1 0 $X=256050 $Y=100160
X9252 1 2 115 504 441 477 123 504 SDFRRQJI3VX1 $T=271600 78400 1 0 $X=271170 $Y=73280
X9253 1 2 123 514 441 477 116 514 SDFRRQJI3VX1 $T=274400 96320 0 0 $X=273970 $Y=95680
X9254 1 2 115 1277 441 514 123 1277 SDFRRQJI3VX1 $T=274960 78400 0 0 $X=274530 $Y=77760
X9255 1 2 111 513 441 514 SPI_CS 513 SDFRRQJI3VX1 $T=274960 87360 1 0 $X=274530 $Y=82240
X9256 1 2 123 527 441 514 116 527 SDFRRQJI3VX1 $T=295120 87360 1 180 $X=274530 $Y=86720
X9257 1 2 713 527 457 911 SPI_CS 911 SDFRRQJI3VX1 $T=274960 132160 1 0 $X=274530 $Y=127040
X9258 1 2 713 477 457 520 SPI_CS 520 SDFRRQJI3VX1 $T=274960 141120 1 0 $X=274530 $Y=136000
X9259 1 2 713 514 457 538 SPI_CS 538 SDFRRQJI3VX1 $T=274960 141120 0 0 $X=274530 $Y=140480
X9260 1 2 113 503 457 524 SPI_CS 503 SDFRRQJI3VX1 $T=295120 150080 0 180 $X=274530 $Y=144960
X9261 1 2 123 519 442 522 116 519 SDFRRQJI3VX1 $T=275520 212800 1 0 $X=275090 $Y=207680
X9262 1 2 123 524 441 526 116 524 SDFRRQJI3VX1 $T=278880 105280 0 0 $X=278450 $Y=104640
X9263 1 2 123 526 441 527 116 526 SDFRRQJI3VX1 $T=278880 114240 1 0 $X=278450 $Y=109120
X9264 1 2 123 522 442 540 116 522 SDFRRQJI3VX1 $T=299040 203840 1 180 $X=278450 $Y=203200
X9265 1 2 1123 925 442 587 98 1123 SDFRRQJI3VX1 $T=310800 185920 0 180 $X=290210 $Y=180800
X9266 1 2 123 535 457 537 116 535 SDFRRQJI3VX1 $T=291760 168000 0 0 $X=291330 $Y=167360
X9267 1 2 123 536 457 535 116 529 SDFRRQJI3VX1 $T=291760 185920 0 0 $X=291330 $Y=185280
X9268 1 2 123 554 457 541 116 540 SDFRRQJI3VX1 $T=312480 203840 0 180 $X=291890 $Y=198720
X9269 1 2 115 558 441 526 123 558 SDFRRQJI3VX1 $T=292880 105280 1 0 $X=292450 $Y=100160
X9270 1 2 123 919 457 529 116 541 SDFRRQJI3VX1 $T=292880 194880 0 0 $X=292450 $Y=194240
X9271 1 2 123 537 457 553 116 537 SDFRRQJI3VX1 $T=314160 114240 1 180 $X=293570 $Y=113600
X9272 1 2 111 1127 441 526 123 1127 SDFRRQJI3VX1 $T=294560 96320 1 0 $X=294130 $Y=91200
X9273 1 2 111 562 441 524 123 562 SDFRRQJI3VX1 $T=295120 87360 1 0 $X=294690 $Y=82240
X9274 1 2 115 563 441 524 123 563 SDFRRQJI3VX1 $T=295120 87360 0 0 $X=294690 $Y=86720
X9275 1 2 123 561 441 524 116 561 SDFRRQJI3VX1 $T=295120 123200 1 0 $X=294690 $Y=118080
X9276 1 2 713 561 457 572 SPI_CS 572 SDFRRQJI3VX1 $T=298480 132160 1 0 $X=298050 $Y=127040
X9277 1 2 713 526 457 573 SPI_CS 573 SDFRRQJI3VX1 $T=298480 141120 1 0 $X=298050 $Y=136000
X9278 1 2 113 565 457 561 SPI_CS 565 SDFRRQJI3VX1 $T=318640 141120 1 180 $X=298050 $Y=140480
X9279 1 2 713 524 457 574 SPI_CS 574 SDFRRQJI3VX1 $T=298480 150080 1 0 $X=298050 $Y=144960
X9280 1 2 123 553 457 669 116 553 SDFRRQJI3VX1 $T=333760 114240 0 180 $X=313170 $Y=109120
X9281 1 2 115 602 457 561 SPI_CS 602 SDFRRQJI3VX1 $T=314720 96320 0 0 $X=314290 $Y=95680
X9282 1 2 123 568 457 561 116 568 SDFRRQJI3VX1 $T=314720 105280 1 0 $X=314290 $Y=100160
X9283 1 2 111 571 457 561 SPI_CS 571 SDFRRQJI3VX1 $T=315840 96320 1 0 $X=315410 $Y=91200
X9284 1 2 113 930 457 568 SPI_CS 930 SDFRRQJI3VX1 $T=316960 114240 0 0 $X=316530 $Y=113600
X9285 1 2 115 606 457 568 SPI_CS 606 SDFRRQJI3VX1 $T=338240 87360 0 180 $X=317650 $Y=82240
X9286 1 2 111 607 457 568 SPI_CS 607 SDFRRQJI3VX1 $T=338800 78400 1 180 $X=318210 $Y=77760
X9287 1 2 111 628 457 626 SPI_CS 628 SDFRRQJI3VX1 $T=351680 69440 1 180 $X=331090 $Y=68800
X9288 1 2 115 629 457 626 SPI_CS 629 SDFRRQJI3VX1 $T=351680 78400 0 180 $X=331090 $Y=73280
X9289 1 2 123 626 457 568 116 626 SDFRRQJI3VX1 $T=352240 87360 1 180 $X=331650 $Y=86720
X9290 1 2 113 597 457 639 SPI_CS 597 SDFRRQJI3VX1 $T=352240 105280 1 180 $X=331650 $Y=104640
X9291 1 2 113 1295 457 626 SPI_CS 1295 SDFRRQJI3VX1 $T=352240 123200 0 180 $X=331650 $Y=118080
X9292 1 2 113 103 457 638 SPI_CS 103 SDFRRQJI3VX1 $T=352240 123200 1 180 $X=331650 $Y=122560
X9293 1 2 115 1157 105 638 SPI_CS 1157 SDFRRQJI3VX1 $T=360080 69440 0 0 $X=359650 $Y=68800
X9294 1 2 111 655 105 638 SPI_CS 655 SDFRRQJI3VX1 $T=360080 78400 1 0 $X=359650 $Y=73280
X9295 1 2 115 952 105 639 SPI_CS 952 SDFRRQJI3VX1 $T=360080 78400 0 0 $X=359650 $Y=77760
X9296 1 2 111 635 105 639 SPI_CS 635 SDFRRQJI3VX1 $T=360080 87360 1 0 $X=359650 $Y=82240
X9297 1 2 123 639 105 626 116 639 SDFRRQJI3VX1 $T=360080 87360 0 0 $X=359650 $Y=86720
X9298 1 2 123 640 105 638 116 640 SDFRRQJI3VX1 $T=360080 96320 1 0 $X=359650 $Y=91200
X9299 1 2 123 638 105 639 116 638 SDFRRQJI3VX1 $T=360080 96320 0 0 $X=359650 $Y=95680
X9300 1 2 113 656 105 637 SPI_CS 656 SDFRRQJI3VX1 $T=360080 114240 0 0 $X=359650 $Y=113600
X9301 1 2 113 657 105 640 SPI_CS 657 SDFRRQJI3VX1 $T=360080 123200 1 0 $X=359650 $Y=118080
X9302 1 2 113 1308 105 633 SPI_CS 1308 SDFRRQJI3VX1 $T=360080 123200 0 0 $X=359650 $Y=122560
X9303 1 2 113 1158 105 669 SPI_CS 1158 SDFRRQJI3VX1 $T=360080 132160 1 0 $X=359650 $Y=127040
X9304 1 2 123 637 105 640 116 637 SDFRRQJI3VX1 $T=361200 105280 1 0 $X=360770 $Y=100160
X9305 1 2 123 633 105 637 116 633 SDFRRQJI3VX1 $T=381360 105280 1 180 $X=360770 $Y=104640
X9306 1 2 123 669 105 633 116 669 SDFRRQJI3VX1 $T=381360 114240 0 180 $X=360770 $Y=109120
X9307 1 2 111 958 105 669 SPI_CS 958 SDFRRQJI3VX1 $T=380240 78400 0 0 $X=379810 $Y=77760
X9308 1 2 115 735 105 669 SPI_CS 735 SDFRRQJI3VX1 $T=380240 87360 1 0 $X=379810 $Y=82240
X9309 1 2 115 736 105 640 SPI_CS 736 SDFRRQJI3VX1 $T=380240 87360 0 0 $X=379810 $Y=86720
X9310 1 2 111 666 105 640 SPI_CS 666 SDFRRQJI3VX1 $T=380240 96320 0 0 $X=379810 $Y=95680
X9311 1 2 696 688 105 687 102 687 SDFRRQJI3VX1 $T=391440 132160 0 0 $X=391010 $Y=131520
X9312 1 2 115 106 105 633 SPI_CS 106 SDFRRQJI3VX1 $T=395360 78400 1 0 $X=394930 $Y=73280
X9313 1 2 115 692 105 637 SPI_CS 692 SDFRRQJI3VX1 $T=395360 96320 1 0 $X=394930 $Y=91200
X9314 1 2 111 1167 105 633 SPI_CS 1167 SDFRRQJI3VX1 $T=400400 87360 1 0 $X=399970 $Y=82240
X9315 1 2 111 107 105 637 SPI_CS 107 SDFRRQJI3VX1 $T=400400 87360 0 0 $X=399970 $Y=86720
X9316 1 2 986 1171 161 NO2JI3VX0 $T=40880 168000 1 180 $X=38210 $Y=167360
X9317 1 2 985 211 751 NO2JI3VX0 $T=44800 159040 0 0 $X=44370 $Y=158400
X9318 1 2 151 176 752 NO2JI3VX0 $T=47040 159040 1 0 $X=46610 $Y=153920
X9319 1 2 991 175 746 NO2JI3VX0 $T=53200 168000 1 180 $X=50530 $Y=167360
X9320 1 2 707 992 1182 NO2JI3VX0 $T=52640 176960 0 0 $X=52210 $Y=176320
X9321 1 2 175 179 992 NO2JI3VX0 $T=53760 168000 1 0 $X=53330 $Y=162880
X9322 1 2 199 1186 192 NO2JI3VX0 $T=62720 185920 0 180 $X=60050 $Y=180800
X9323 1 2 167 764 201 NO2JI3VX0 $T=62160 159040 1 0 $X=61730 $Y=153920
X9324 1 2 210 767 215 NO2JI3VX0 $T=69440 185920 0 180 $X=66770 $Y=180800
X9325 1 2 210 999 203 NO2JI3VX0 $T=71680 203840 0 180 $X=69010 $Y=198720
X9326 1 2 178 1195 212 NO2JI3VX0 $T=77840 194880 1 0 $X=77410 $Y=189760
X9327 1 2 1195 219 220 NO2JI3VX0 $T=80640 185920 1 180 $X=77970 $Y=185280
X9328 1 2 810 1038 825 NO2JI3VX0 $T=148960 123200 1 0 $X=148530 $Y=118080
X9329 1 2 343 1377 1058 NO2JI3VX0 $T=179200 176960 1 180 $X=176530 $Y=176320
X9330 1 2 842 378 361 NO2JI3VX0 $T=179760 203840 1 0 $X=179330 $Y=198720
X9331 1 2 1411 1065 122 NO2JI3VX0 $T=184800 185920 1 0 $X=184370 $Y=180800
X9332 1 2 839 400 856 NO2JI3VX0 $T=204960 185920 1 180 $X=202290 $Y=185280
X9333 1 2 133 1392 859 NO2JI3VX0 $T=218960 176960 0 180 $X=216290 $Y=171840
X9334 1 2 720 421 97 NO2JI3VX0 $T=220080 185920 0 180 $X=217410 $Y=180800
X9335 1 2 883 1098 446 NO2JI3VX0 $T=239680 168000 1 0 $X=239250 $Y=162880
X9336 1 2 135 1100 1256 NO2JI3VX0 $T=240240 194880 0 0 $X=239810 $Y=194240
X9337 1 2 485 135 440 NO2JI3VX0 $T=244720 194880 1 180 $X=242050 $Y=194240
X9338 1 2 1093 890 883 NO2JI3VX0 $T=245280 176960 0 180 $X=242610 $Y=171840
X9339 1 2 893 466 459 NO2JI3VX0 $T=253120 176960 1 180 $X=250450 $Y=176320
X9340 1 2 1258 463 893 NO2JI3VX0 $T=253120 185920 0 180 $X=250450 $Y=180800
X9341 1 2 472 1109 895 NO2JI3VX0 $T=255360 168000 0 0 $X=254930 $Y=167360
X9342 1 2 1111 478 476 NO2JI3VX0 $T=261520 185920 0 180 $X=258850 $Y=180800
X9343 1 2 584 933 588 NO2JI3VX0 $T=324800 24640 1 0 $X=324370 $Y=19520
X9344 1 2 1410 1351 1298 NO2JI3VX0 $T=330960 168000 1 180 $X=328290 $Y=167360
X9345 1 2 612 939 617 NO2JI3VX0 $T=337680 159040 1 0 $X=337250 $Y=153920
X9346 1 2 917 614 605 NO2JI3VX0 $T=338800 24640 0 0 $X=338370 $Y=24000
X9347 1 2 1402 1353 613 NO2JI3VX0 $T=339360 212800 0 0 $X=338930 $Y=212160
X9348 1 2 946 945 612 NO2JI3VX0 $T=343840 176960 1 180 $X=341170 $Y=176320
X9349 1 2 622 613 1389 NO2JI3VX0 $T=349440 212800 1 180 $X=346770 $Y=212160
X9350 1 2 627 1175 950 NO2JI3VX0 $T=352240 159040 1 180 $X=349570 $Y=158400
X9351 1 2 652 141 658 NO2JI3VX0 $T=380240 24640 0 180 $X=377570 $Y=19520
X9352 1 2 672 1386 681 NO2JI3VX0 $T=384720 114240 0 0 $X=384290 $Y=113600
X9353 1 2 679 1365 674 NO2JI3VX0 $T=384720 141120 0 0 $X=384290 $Y=140480
X9354 1 2 671 1358 609 NO2JI3VX0 $T=385280 159040 1 0 $X=384850 $Y=153920
X9355 1 2 675 672 687 NO2JI3VX0 $T=392000 105280 1 180 $X=389330 $Y=104640
X9356 1 2 697 949 1160 NO2JI3VX0 $T=393680 24640 0 180 $X=391010 $Y=19520
X9357 1 2 85 110 755 995 1180 NA4JI3VX0 $T=54320 159040 1 180 $X=49970 $Y=158400
X9358 1 2 1412 855 391 399 853 NA4JI3VX0 $T=198240 185920 1 0 $X=197810 $Y=180800
X9359 1 2 949 621 614 933 141 NA4JI3VX0 $T=347760 24640 1 0 $X=347330 $Y=19520
X9360 1 2 1161 1413 682 677 680 NA4JI3VX0 $T=394240 141120 0 180 $X=389890 $Y=136000
X9361 1 2 157 1414 150 NA2JI3VX0 $T=26320 168000 1 0 $X=25890 $Y=162880
X9362 1 2 165 1406 1176 NA2JI3VX0 $T=33600 150080 0 0 $X=33170 $Y=149440
X9363 1 2 157 1407 169 NA2JI3VX0 $T=42000 176960 1 180 $X=39330 $Y=176320
X9364 1 2 747 989 988 NA2JI3VX0 $T=40880 159040 0 0 $X=40450 $Y=158400
X9365 1 2 1369 168 1177 NA2JI3VX0 $T=42000 150080 0 0 $X=41570 $Y=149440
X9366 1 2 752 755 151 NA2JI3VX0 $T=49840 150080 1 180 $X=47170 $Y=149440
X9367 1 2 751 995 985 NA2JI3VX0 $T=47600 159040 0 0 $X=47170 $Y=158400
X9368 1 2 753 706 1186 NA2JI3VX0 $T=52080 185920 1 0 $X=51650 $Y=180800
X9369 1 2 992 758 174 NA2JI3VX0 $T=53760 176960 1 0 $X=53330 $Y=171840
X9370 1 2 201 766 167 NA2JI3VX0 $T=67760 159040 0 180 $X=65090 $Y=153920
X9371 1 2 1394 998 1188 NA2JI3VX0 $T=71120 168000 1 180 $X=68450 $Y=167360
X9372 1 2 236 226 227 NA2JI3VX0 $T=90160 24640 1 180 $X=87490 $Y=24000
X9373 1 2 773 1341 227 NA2JI3VX0 $T=91280 42560 0 180 $X=88610 $Y=37440
X9374 1 2 232 228 227 NA2JI3VX0 $T=92400 42560 1 0 $X=91970 $Y=37440
X9375 1 2 776 784 227 NA2JI3VX0 $T=103600 24640 0 0 $X=103170 $Y=24000
X9376 1 2 242 787 227 NA2JI3VX0 $T=110320 24640 1 180 $X=107650 $Y=24000
X9377 1 2 252 796 227 NA2JI3VX0 $T=115360 24640 1 180 $X=112690 $Y=24000
X9378 1 2 268 1207 227 NA2JI3VX0 $T=124880 33600 1 0 $X=124450 $Y=28480
X9379 1 2 279 805 227 NA2JI3VX0 $T=135520 33600 1 180 $X=132850 $Y=32960
X9380 1 2 284 1020 286 NA2JI3VX0 $T=133280 114240 0 0 $X=132850 $Y=113600
X9381 1 2 273 295 286 NA2JI3VX0 $T=143920 114240 0 0 $X=143490 $Y=113600
X9382 1 2 299 297 227 NA2JI3VX0 $T=147840 24640 1 180 $X=145170 $Y=24000
X9383 1 2 1218 90 549 NA2JI3VX0 $T=148400 114240 1 180 $X=145730 $Y=113600
X9384 1 2 1361 300 549 NA2JI3VX0 $T=148960 123200 0 180 $X=146290 $Y=118080
X9385 1 2 812 818 227 NA2JI3VX0 $T=148960 33600 0 0 $X=148530 $Y=32960
X9386 1 2 1033 1037 286 NA2JI3VX0 $T=148960 114240 1 0 $X=148530 $Y=109120
X9387 1 2 1026 120 286 NA2JI3VX0 $T=152320 105280 0 0 $X=151890 $Y=104640
X9388 1 2 323 1173 227 NA2JI3VX0 $T=160720 33600 0 180 $X=158050 $Y=28480
X9389 1 2 1047 1044 549 NA2JI3VX0 $T=161840 114240 0 180 $X=159170 $Y=109120
X9390 1 2 1004 1322 286 NA2JI3VX0 $T=164640 114240 1 0 $X=164210 $Y=109120
X9391 1 2 342 1321 227 NA2JI3VX0 $T=170240 33600 1 0 $X=169810 $Y=28480
X9392 1 2 356 1230 286 NA2JI3VX0 $T=175840 123200 1 0 $X=175410 $Y=118080
X9393 1 2 364 360 362 NA2JI3VX0 $T=183680 194880 0 180 $X=181010 $Y=189760
X9394 1 2 365 363 227 NA2JI3VX0 $T=182560 33600 0 0 $X=182130 $Y=32960
X9395 1 2 839 1344 1415 NA2JI3VX0 $T=183120 176960 1 0 $X=182690 $Y=171840
X9396 1 2 407 846 1415 NA2JI3VX0 $T=189280 176960 0 180 $X=186610 $Y=171840
X9397 1 2 847 376 369 NA2JI3VX0 $T=189840 194880 1 180 $X=187170 $Y=194240
X9398 1 2 384 382 1379 NA2JI3VX0 $T=195440 176960 1 0 $X=195010 $Y=171840
X9399 1 2 856 1236 839 NA2JI3VX0 $T=202160 185920 1 180 $X=199490 $Y=185280
X9400 1 2 402 393 227 NA2JI3VX0 $T=203280 42560 1 180 $X=200610 $Y=41920
X9401 1 2 395 416 128 NA2JI3VX0 $T=206080 203840 0 0 $X=205650 $Y=203200
X9402 1 2 862 411 227 NA2JI3VX0 $T=211120 33600 1 180 $X=208450 $Y=32960
X9403 1 2 127 1416 425 NA2JI3VX0 $T=211120 185920 0 180 $X=208450 $Y=180800
X9404 1 2 reset_l 1409 865 NA2JI3VX0 $T=211680 212800 0 0 $X=211250 $Y=212160
X9405 1 2 1080 1248 1084 NA2JI3VX0 $T=212800 203840 1 0 $X=212370 $Y=198720
X9406 1 2 444 866 447 NA2JI3VX0 $T=213920 33600 0 0 $X=213490 $Y=32960
X9407 1 2 97 425 1392 NA2JI3VX0 $T=216720 176960 0 180 $X=214050 $Y=171840
X9408 1 2 127 414 421 NA2JI3VX0 $T=220080 159040 1 0 $X=219650 $Y=153920
X9409 1 2 1096 880 447 NA2JI3VX0 $T=235760 33600 0 180 $X=233090 $Y=28480
X9410 1 2 1090 1250 1084 NA2JI3VX0 $T=237440 203840 0 180 $X=234770 $Y=198720
X9411 1 2 881 1349 447 NA2JI3VX0 $T=244160 33600 0 180 $X=241490 $Y=28480
X9412 1 2 1103 889 448 NA2JI3VX0 $T=248080 168000 1 180 $X=245410 $Y=167360
X9413 1 2 888 1258 890 NA2JI3VX0 $T=248640 185920 0 180 $X=245970 $Y=180800
X9414 1 2 461 1334 447 NA2JI3VX0 $T=253120 33600 0 0 $X=252690 $Y=32960
X9415 1 2 1096 897 521 NA2JI3VX0 $T=257040 42560 1 0 $X=256610 $Y=37440
X9416 1 2 475 1350 447 NA2JI3VX0 $T=261520 33600 1 0 $X=261090 $Y=28480
X9417 1 2 493 902 492 NA2JI3VX0 $T=269920 185920 1 180 $X=267250 $Y=185280
X9418 1 2 100 903 483 NA2JI3VX0 $T=268800 194880 1 0 $X=268370 $Y=189760
X9419 1 2 1381 906 904 NA2JI3VX0 $T=270480 176960 0 0 $X=270050 $Y=176320
X9420 1 2 501 907 447 NA2JI3VX0 $T=272160 42560 1 0 $X=271730 $Y=37440
X9421 1 2 515 511 508 NA2JI3VX0 $T=277760 185920 0 180 $X=275090 $Y=180800
X9422 1 2 506 910 508 NA2JI3VX0 $T=275520 185920 0 0 $X=275090 $Y=185280
X9423 1 2 516 500 447 NA2JI3VX0 $T=278320 33600 0 180 $X=275650 $Y=28480
X9424 1 2 517 901 447 NA2JI3VX0 $T=278320 42560 0 180 $X=275650 $Y=37440
X9425 1 2 512 913 447 NA2JI3VX0 $T=278320 24640 0 0 $X=277890 $Y=24000
X9426 1 2 127 1244 539 NA2JI3VX0 $T=281120 168000 0 0 $X=280690 $Y=167360
X9427 1 2 517 914 521 NA2JI3VX0 $T=282240 42560 1 0 $X=281810 $Y=37440
X9428 1 2 516 528 521 NA2JI3VX0 $T=282800 33600 1 0 $X=282370 $Y=28480
X9429 1 2 531 1280 447 NA2JI3VX0 $T=295680 24640 1 180 $X=293010 $Y=24000
X9430 1 2 1125 1281 447 NA2JI3VX0 $T=295680 33600 1 180 $X=293010 $Y=32960
X9431 1 2 127 1417 544 NA2JI3VX0 $T=297920 176960 1 0 $X=297490 $Y=171840
X9432 1 2 553 543 542 NA2JI3VX0 $T=302960 123200 0 0 $X=302530 $Y=122560
X9433 1 2 570 926 447 NA2JI3VX0 $T=313040 33600 1 180 $X=310370 $Y=32960
X9434 1 2 559 546 566 NA2JI3VX0 $T=313040 212800 0 0 $X=312610 $Y=212160
X9435 1 2 560 929 447 NA2JI3VX0 $T=316960 33600 1 0 $X=316530 $Y=28480
X9436 1 2 585 582 931 NA2JI3VX0 $T=321440 168000 1 0 $X=321010 $Y=162880
X9437 1 2 591 601 1297 NA2JI3VX0 $T=329840 176960 0 0 $X=329410 $Y=176320
X9438 1 2 600 938 598 NA2JI3VX0 $T=330960 194880 1 0 $X=330530 $Y=189760
X9439 1 2 592 936 447 NA2JI3VX0 $T=332080 33600 0 0 $X=331650 $Y=32960
X9440 1 2 594 1303 447 NA2JI3VX0 $T=337120 33600 1 0 $X=336690 $Y=28480
X9441 1 2 592 138 521 NA2JI3VX0 $T=337120 42560 1 0 $X=336690 $Y=37440
X9442 1 2 616 1384 521 NA2JI3VX0 $T=343280 42560 1 0 $X=342850 $Y=37440
X9443 1 2 616 1307 447 NA2JI3VX0 $T=345520 42560 1 0 $X=345090 $Y=37440
X9444 1 2 1149 951 447 NA2JI3VX0 $T=349440 51520 1 0 $X=349010 $Y=46400
X9445 1 2 950 623 627 NA2JI3VX0 $T=351680 168000 0 180 $X=349010 $Y=162880
X9446 1 2 642 943 1146 NA2JI3VX0 $T=365680 176960 0 180 $X=363010 $Y=171840
X9447 1 2 636 641 643 NA2JI3VX0 $T=363440 185920 1 0 $X=363010 $Y=180800
X9448 1 2 954 142 643 NA2JI3VX0 $T=367920 185920 0 180 $X=365250 $Y=180800
X9449 1 2 732 1354 447 NA2JI3VX0 $T=366240 42560 1 0 $X=365810 $Y=37440
X9450 1 2 143 1355 447 NA2JI3VX0 $T=370720 42560 0 180 $X=368050 $Y=37440
X9451 1 2 732 1356 521 NA2JI3VX0 $T=372960 42560 0 180 $X=370290 $Y=37440
X9452 1 2 645 1152 447 NA2JI3VX0 $T=371840 33600 1 0 $X=371410 $Y=28480
X9453 1 2 653 1364 447 NA2JI3VX0 $T=375200 42560 0 180 $X=372530 $Y=37440
X9454 1 2 653 1156 521 NA2JI3VX0 $T=376880 42560 1 0 $X=376450 $Y=37440
X9455 1 2 650 1339 447 NA2JI3VX0 $T=377440 33600 0 0 $X=377010 $Y=32960
X9456 1 2 661 665 1385 NA2JI3VX0 $T=385840 159040 1 180 $X=383170 $Y=158400
X9457 1 2 681 1408 676 NA2JI3VX0 $T=385840 123200 1 0 $X=385410 $Y=118080
X9458 1 2 673 677 661 NA2JI3VX0 $T=389200 141120 0 180 $X=386530 $Y=136000
X9459 1 2 689 1162 447 NA2JI3VX0 $T=396480 33600 0 180 $X=393810 $Y=28480
X9460 1 2 691 962 447 NA2JI3VX0 $T=396480 33600 1 180 $X=393810 $Y=32960
X9461 1 2 662 682 966 NA2JI3VX0 $T=395360 150080 1 0 $X=394930 $Y=144960
X9462 1 2 1159 967 1165 NA2JI3VX0 $T=395920 159040 0 0 $X=395490 $Y=158400
X9463 1 2 1166 696 1413 NA2JI3VX0 $T=402080 141120 0 180 $X=399410 $Y=136000
X9464 1 2 1418 716 228 down_switches<4> ON21JI3VX4 $T=91280 42560 1 180 $X=82450 $Y=41920
X9465 1 2 114 716 226 down_switches<1> ON21JI3VX4 $T=84560 24640 1 0 $X=84130 $Y=19520
X9466 1 2 1419 716 1341 down_switches<2> ON21JI3VX4 $T=87360 33600 0 0 $X=86930 $Y=32960
X9467 1 2 1006 716 784 down_switches<3> ON21JI3VX4 $T=109760 24640 0 180 $X=100930 $Y=19520
X9468 1 2 786 716 787 down_switches<5> ON21JI3VX4 $T=109760 24640 1 0 $X=109330 $Y=19520
X9469 1 2 793 716 796 down_switches<6> ON21JI3VX4 $T=118160 24640 1 0 $X=117730 $Y=19520
X9470 1 2 1015 716 1207 down_switches<7> ON21JI3VX4 $T=134960 24640 0 180 $X=126130 $Y=19520
X9471 1 2 809 716 805 down_switches<9> ON21JI3VX4 $T=137200 33600 0 180 $X=128370 $Y=28480
X9472 1 2 1420 716 297 down_switches<8> ON21JI3VX4 $T=140000 24640 1 180 $X=131170 $Y=24000
X9473 1 2 314 716 818 down_switches<0> ON21JI3VX4 $T=154560 33600 0 180 $X=145730 $Y=28480
X9474 1 2 1421 716 1173 down_switches<10> ON21JI3VX4 $T=160720 24640 0 180 $X=151890 $Y=19520
X9475 1 2 341 716 1321 down_switches<11> ON21JI3VX4 $T=170240 24640 1 180 $X=161410 $Y=24000
X9476 1 2 1422 716 363 down_switches<12> ON21JI3VX4 $T=183120 33600 0 180 $X=174290 $Y=28480
X9477 1 2 412 716 393 down_switches<13> ON21JI3VX4 $T=201600 42560 0 180 $X=192770 $Y=37440
X9478 1 2 1077 716 411 down_switches<14> ON21JI3VX4 $T=207760 33600 0 180 $X=198930 $Y=28480
X9479 1 2 1423 716 866 down_switches<15> ON21JI3VX4 $T=218960 33600 0 180 $X=210130 $Y=28480
X9480 1 2 1330 716 880 down_switches<17> ON21JI3VX4 $T=239120 24640 0 180 $X=230290 $Y=19520
X9481 1 2 1424 716 1349 down_switches<16> ON21JI3VX4 $T=241360 24640 1 180 $X=232530 $Y=24000
X9482 1 2 1425 716 1350 down_switches<20> ON21JI3VX4 $T=266560 24640 1 180 $X=257730 $Y=24000
X9483 1 2 1118 716 901 down_switches<18> ON21JI3VX4 $T=270480 42560 0 180 $X=261650 $Y=37440
X9484 1 2 1426 716 500 down_switches<19> ON21JI3VX4 $T=274960 33600 1 180 $X=266130 $Y=32960
X9485 1 2 1427 716 1280 down_switches<21> ON21JI3VX4 $T=296240 24640 0 180 $X=287410 $Y=19520
X9486 1 2 1126 716 1281 down_switches<22> ON21JI3VX4 $T=296240 33600 0 180 $X=287410 $Y=28480
X9487 1 2 567 716 926 down_switches<23> ON21JI3VX4 $T=317520 24640 1 180 $X=308690 $Y=24000
X9488 1 2 1133 716 929 down_switches<24> ON21JI3VX4 $T=322000 24640 0 180 $X=313170 $Y=19520
X9489 1 2 937 716 936 down_switches<25> ON21JI3VX4 $T=337120 24640 1 180 $X=328290 $Y=24000
X9490 1 2 624 716 1307 down_switches<26> ON21JI3VX4 $T=351120 33600 1 180 $X=342290 $Y=32960
X9491 1 2 1428 716 1354 down_switches<27> ON21JI3VX4 $T=366240 33600 1 180 $X=357410 $Y=32960
X9492 1 2 1309 716 1364 down_switches<28> ON21JI3VX4 $T=366240 42560 0 180 $X=357410 $Y=37440
X9493 1 2 648 716 1152 down_switches<31> ON21JI3VX4 $T=376880 24640 0 180 $X=368050 $Y=19520
X9494 1 2 684 716 962 down_switches<30> ON21JI3VX4 $T=393680 33600 1 180 $X=384850 $Y=32960
X9495 1 2 1429 716 1162 down_switches<29> ON21JI3VX4 $T=386960 24640 0 0 $X=386530 $Y=24000
X9496 1 2 196 284 1366 AND2JI3VX1 $T=61600 33600 1 0 $X=61170 $Y=28480
X9497 1 2 196 273 206 AND2JI3VX1 $T=62160 24640 0 0 $X=61730 $Y=24000
X9498 1 2 196 1004 1367 AND2JI3VX1 $T=75600 33600 1 0 $X=75170 $Y=28480
X9499 1 2 196 1026 777 AND2JI3VX1 $T=137760 33600 1 0 $X=137330 $Y=28480
X9500 1 2 196 1033 778 AND2JI3VX1 $T=142240 24640 0 0 $X=141810 $Y=24000
X9501 1 2 196 356 357 AND2JI3VX1 $T=180320 24640 1 180 $X=176530 $Y=24000
X9502 1 2 410 978 545 548 615 NA4JI3VX2 $T=306320 24640 1 180 $X=298610 $Y=24000
X9503 1 2 521 488 447 NO2I1JI3VX2 $T=313040 33600 0 180 $X=307570 $Y=28480
X9504 1 2 1038 1216 290 EO2JI3VX0 $T=141680 123200 0 180 $X=135650 $Y=118080
X9505 1 2 1391 312 1430 EO2JI3VX0 $T=156240 132160 0 180 $X=150210 $Y=127040
X9506 1 2 364 362 1403 EO2JI3VX0 $T=181440 194880 0 180 $X=175410 $Y=189760
X9507 1 2 395 128 1404 EO2JI3VX0 $T=194320 203840 0 0 $X=193890 $Y=203200
X9508 1 2 100 483 507 EO2JI3VX0 $T=271040 203840 1 0 $X=270610 $Y=198720
X9509 1 2 519 IC_addr<1> 534 EO2JI3VX0 $T=278880 212800 0 0 $X=278450 $Y=212160
X9510 1 2 522 IC_addr<0> 1398 EO2JI3VX0 $T=286720 212800 0 0 $X=286290 $Y=212160
X9511 1 2 591 1297 579 EO2JI3VX0 $T=328160 176960 0 180 $X=322130 $Y=171840
X9512 1 2 161 745 172 AND2JI3VX0 $T=41440 168000 0 0 $X=41010 $Y=167360
X9513 1 2 186 766 1180 AND2JI3VX0 $T=61600 159040 0 180 $X=57810 $Y=153920
X9514 1 2 129 1286 1247 AND2JI3VX0 $T=211680 168000 1 0 $X=211250 $Y=162880
X9515 1 2 893 459 452 AND2JI3VX0 $T=250320 176960 1 180 $X=246530 $Y=176320
X9516 1 2 463 456 1401 AND2JI3VX0 $T=250880 194880 0 0 $X=250450 $Y=194240
X9517 1 2 521 881 1261 AND2JI3VX0 $T=255920 33600 0 180 $X=252130 $Y=28480
X9518 1 2 622 730 1402 AND2JI3VX0 $T=346640 212800 1 180 $X=342850 $Y=212160
X9519 1 2 521 645 663 AND2JI3VX0 $T=384160 33600 0 180 $X=380370 $Y=28480
X9520 1 2 960 677 671 AND2JI3VX0 $T=389200 150080 0 180 $X=385410 $Y=144960
X9521 1 2 521 689 968 AND2JI3VX0 $T=397040 33600 1 0 $X=396610 $Y=28480
X9522 1 2 521 691 973 AND2JI3VX0 $T=400400 33600 0 0 $X=399970 $Y=32960
X9523 1 2 707 1186 1184 192 753 AN22JI3VX1 $T=59360 185920 0 180 $X=55010 $Y=180800
X9524 1 2 212 999 205 210 203 AN22JI3VX1 $T=71680 194880 1 180 $X=67330 $Y=194240
X9525 1 2 215 210 996 214 213 AN22JI3VX1 $T=74480 176960 1 180 $X=70130 $Y=176320
X9526 1 2 290 304 1375 418 1017 AN22JI3VX1 $T=137200 114240 0 0 $X=136770 $Y=113600
X9527 1 2 1210 304 1025 418 1019 AN22JI3VX1 $T=142240 132160 0 180 $X=137890 $Y=127040
X9528 1 2 1430 304 119 418 296 AN22JI3VX1 $T=150080 132160 0 180 $X=145730 $Y=127040
X9529 1 2 367 549 1043 418 309 AN22JI3VX1 $T=154560 123200 1 0 $X=154130 $Y=118080
X9530 1 2 348 549 344 418 335 AN22JI3VX1 $T=172480 132160 0 180 $X=168130 $Y=127040
X9531 1 2 373 549 1061 418 349 AN22JI3VX1 $T=184240 132160 0 180 $X=179890 $Y=127040
X9532 1 2 368 844 1068 842 361 AN22JI3VX1 $T=187040 203840 0 180 $X=182690 $Y=198720
X9533 1 2 862 318 545 227 413 AN22JI3VX1 $T=223440 33600 1 180 $X=219090 $Y=32960
X9534 1 2 856 1080 873 132 453 AN22JI3VX1 $T=223440 185920 1 180 $X=219090 $Y=185280
X9535 1 2 444 318 548 447 428 AN22JI3VX1 $T=240800 33600 0 180 $X=236450 $Y=28480
X9536 1 2 446 883 467 1093 886 AN22JI3VX1 $T=238000 159040 0 0 $X=237570 $Y=158400
X9537 1 2 448 890 1331 883 888 AN22JI3VX1 $T=241920 176960 0 0 $X=241490 $Y=176320
X9538 1 2 472 463 462 456 893 AN22JI3VX1 $T=254240 185920 1 180 $X=249890 $Y=185280
X9539 1 2 1125 488 978 447 920 AN22JI3VX1 $T=297920 33600 0 0 $X=297490 $Y=32960
X9540 1 2 1139 1138 927 603 943 AN22JI3VX1 $T=344960 168000 1 180 $X=340610 $Y=167360
X9541 1 2 659 664 961 668 674 AN22JI3VX1 $T=380240 132160 0 0 $X=379810 $Y=131520
X9542 1 2 659 667 680 679 674 AN22JI3VX1 $T=383040 141120 1 0 $X=382610 $Y=136000
X9543 1 2 678 961 675 670 673 AN22JI3VX1 $T=389760 123200 1 180 $X=385410 $Y=122560
X9544 1 2 537 543 713 NO2JI3VX2 $T=301280 123200 1 180 $X=296370 $Y=122560
X9545 1 2 220 212 1195 1005 AO21JI3VX1 $T=80640 194880 1 0 $X=80210 $Y=189760
X9546 1 2 825 810 1038 1210 AO21JI3VX1 $T=146720 123200 0 180 $X=141810 $Y=118080
X9547 1 2 1431 1058 390 1388 AO21JI3VX1 $T=186480 176960 0 0 $X=186050 $Y=176320
X9548 1 2 440 1256 135 436 AO21JI3VX1 $T=240240 194880 1 180 $X=235330 $Y=194240
X9549 1 2 601 587 925 598 AO21JI3VX1 $T=327040 185920 1 0 $X=326610 $Y=180800
X9550 1 2 623 939 1175 1139 AO21JI3VX1 $T=348320 159040 1 180 $X=343410 $Y=158400
X9551 1 2 947 587 925 643 AO21JI3VX1 $T=345520 185920 1 0 $X=345090 $Y=180800
X9552 1 2 447 671 609 959 AO21JI3VX1 $T=375760 159040 1 0 $X=375330 $Y=153920
X9553 1 2 543 115 537 NA2I1JI3VX2 $T=300720 105280 0 0 $X=300290 $Y=104640
X9554 1 2 537 113 1130 NA2I1JI3VX2 $T=313040 123200 0 0 $X=312610 $Y=122560
X9555 1 2 986 152 enable 169 NA22JI3VX1 $T=40880 176960 1 0 $X=40450 $Y=171840
X9556 1 2 192 759 174 760 NA22JI3VX1 $T=61040 176960 0 180 $X=56690 $Y=171840
X9557 1 2 360 313 382 1415 NA22JI3VX1 $T=179200 176960 1 0 $X=178770 $Y=171840
X9558 1 2 416 319 718 1084 NA22JI3VX1 $T=204400 203840 1 0 $X=203970 $Y=198720
X9559 1 2 476 1111 473 470 NA22JI3VX1 $T=258720 176960 1 180 $X=254370 $Y=176320
X9560 1 2 903 1170 906 508 NA22JI3VX1 $T=271040 185920 0 0 $X=270610 $Y=185280
X9561 1 2 1142 104 943 140 NA22JI3VX1 $T=348880 168000 0 0 $X=348450 $Y=167360
X9562 1 2 675 690 1166 108 NA22JI3VX1 $T=394800 105280 0 0 $X=394370 $Y=104640
X9563 1 2 447 1261 471 588 MU2JI3VX0 $T=250320 24640 0 0 $X=249890 $Y=24000
X9564 1 2 447 663 647 697 MU2JI3VX0 $T=380240 24640 0 0 $X=379810 $Y=24000
X9565 1 2 447 968 694 652 MU2JI3VX0 $T=402640 24640 1 180 $X=396610 $Y=24000
X9566 1 2 447 973 971 1160 MU2JI3VX0 $T=408240 33600 0 180 $X=402210 $Y=28480
X9567 1 2 374 429 221 381 OR3JI3VX1 $T=188160 33600 1 0 $X=187730 $Y=28480
X9568 1 2 401 1346 848 857 OR3JI3VX1 $T=202720 194880 1 0 $X=202290 $Y=189760
X9569 1 2 498 478 1109 899 OR3JI3VX1 $T=258720 168000 0 0 $X=258290 $Y=167360
X9570 1 2 899 1393 898 1432 OR3JI3VX1 $T=263200 168000 0 180 $X=258850 $Y=162880
X9571 1 2 924 632 934 1140 OR3JI3VX1 $T=350000 33600 0 180 $X=345650 $Y=28480
X9572 1 2 211 757 176 1180 755 ON211JI3VX1 $T=49840 159040 1 0 $X=49410 $Y=153920
X9573 1 2 172 85 1315 1317 758 ON211JI3VX1 $T=54320 168000 0 0 $X=53890 $Y=167360
X9574 1 2 213 1397 214 1191 998 ON211JI3VX1 $T=72800 176960 0 180 $X=68450 $Y=171840
X9575 1 2 315 1042 351 1037 1043 ON211JI3VX1 $T=154000 114240 1 0 $X=153570 $Y=109120
X9576 1 2 351 831 833 1322 344 ON211JI3VX1 $T=166880 114240 0 0 $X=166450 $Y=113600
X9577 1 2 351 843 832 1230 1061 ON211JI3VX1 $T=178080 123200 1 0 $X=177650 $Y=118080
X9578 1 2 847 848 369 94 849 ON211JI3VX1 $T=190960 194880 0 0 $X=190530 $Y=194240
X9579 1 2 376 850 378 1068 852 ON211JI3VX1 $T=191520 203840 1 0 $X=191090 $Y=198720
X9580 1 2 1243 130 849 850 1073 ON211JI3VX1 $T=196000 194880 0 0 $X=195570 $Y=194240
X9581 1 2 390 384 124 421 399 ON211JI3VX1 $T=198800 176960 0 0 $X=198370 $Y=176320
X9582 1 2 414 1363 855 1246 1247 ON211JI3VX1 $T=207200 168000 1 0 $X=206770 $Y=162880
X9583 1 2 127 1433 420 1085 1434 ON211JI3VX1 $T=218960 159040 0 180 $X=214610 $Y=153920
X9584 1 2 220 1251 1348 1085 414 ON211JI3VX1 $T=220640 168000 0 180 $X=216290 $Y=162880
X9585 1 2 905 904 1272 1116 495 ON211JI3VX1 $T=273280 176960 0 180 $X=268930 $Y=171840
X9586 1 2 674 678 668 1312 662 ON211JI3VX1 $T=385840 132160 1 0 $X=385410 $Y=127040
X9587 1 2 1414 152 983 169 AN21JI3VX1 $T=29680 168000 1 0 $X=29250 $Y=162880
X9588 1 2 175 989 1315 750 AN21JI3VX1 $T=49840 168000 1 0 $X=49410 $Y=162880
X9589 1 2 1182 707 761 760 AN21JI3VX1 $T=56560 176960 0 0 $X=56130 $Y=176320
X9590 1 2 199 152 1390 220 AN21JI3VX1 $T=66640 185920 1 180 $X=62850 $Y=185280
X9591 1 2 1342 1035 312 303 AN21JI3VX1 $T=150080 123200 0 0 $X=149650 $Y=122560
X9592 1 2 91 1221 824 320 AN21JI3VX1 $T=154560 123200 0 0 $X=154130 $Y=122560
X9593 1 2 840 1232 1411 347 AN21JI3VX1 $T=180880 185920 1 0 $X=180450 $Y=180800
X9594 1 2 839 1060 1378 407 AN21JI3VX1 $T=184800 168000 0 0 $X=184370 $Y=167360
X9595 1 2 847 1238 1069 400 AN21JI3VX1 $T=194320 194880 0 180 $X=190530 $Y=189760
X9596 1 2 1416 1244 125 408 AN21JI3VX1 $T=207200 185920 0 180 $X=203410 $Y=180800
X9597 1 2 1080 130 131 96 AN21JI3VX1 $T=210560 194880 0 0 $X=210130 $Y=194240
X9598 1 2 1116 869 1348 1079 AN21JI3VX1 $T=216160 168000 0 0 $X=215730 $Y=167360
X9599 1 2 1080 1081 1086 1090 AN21JI3VX1 $T=222880 194880 1 180 $X=219090 $Y=194240
X9600 1 2 1258 1170 1263 1256 AN21JI3VX1 $T=245840 194880 0 180 $X=242050 $Y=189760
X9601 1 2 1099 1101 885 452 AN21JI3VX1 $T=243040 168000 1 0 $X=242610 $Y=162880
X9602 1 2 895 472 1105 470 AN21JI3VX1 $T=256480 176960 0 180 $X=252690 $Y=171840
X9603 1 2 1268 1112 473 481 AN21JI3VX1 $T=263200 185920 1 180 $X=259410 $Y=185280
X9604 1 2 1109 1267 1113 1114 AN21JI3VX1 $T=260400 176960 1 0 $X=259970 $Y=171840
X9605 1 2 506 523 1382 515 AN21JI3VX1 $T=281680 185920 0 180 $X=277890 $Y=180800
X9606 1 2 1417 1244 925 136 AN21JI3VX1 $T=302960 176960 1 0 $X=302530 $Y=171840
X9607 1 2 927 557 136 544 AN21JI3VX1 $T=312480 176960 0 180 $X=308690 $Y=171840
X9608 1 2 575 581 1383 599 AN21JI3VX1 $T=322560 168000 1 180 $X=318770 $Y=167360
X9609 1 2 580 1132 935 1175 AN21JI3VX1 $T=338240 159040 0 0 $X=337810 $Y=158400
X9610 1 2 636 1145 1144 954 AN21JI3VX1 $T=362880 176960 1 180 $X=359090 $Y=176320
X9611 1 2 447 671 981 609 AN21JI3VX1 $T=380800 159040 1 0 $X=380370 $Y=153920
X9612 1 2 690 675 145 687 AN21JI3VX1 $T=394240 114240 1 0 $X=393810 $Y=109120
X9613 1 2 150 985 INJI3VX0 $T=33600 168000 1 0 $X=33170 $Y=162880
X9614 1 2 160 151 INJI3VX0 $T=38640 159040 0 180 $X=36530 $Y=153920
X9615 1 2 1171 156 INJI3VX0 $T=38640 168000 1 180 $X=36530 $Y=167360
X9616 1 2 157 161 INJI3VX0 $T=38640 176960 1 0 $X=38210 $Y=171840
X9617 1 2 989 1178 INJI3VX0 $T=47040 168000 1 0 $X=46610 $Y=162880
X9618 1 2 753 707 INJI3VX0 $T=52080 185920 0 0 $X=51650 $Y=185280
X9619 1 2 178 152 INJI3VX0 $T=56560 176960 1 180 $X=54450 $Y=176320
X9620 1 2 194 197 INJI3VX0 $T=63280 150080 1 180 $X=61170 $Y=149440
X9621 1 2 203 1188 INJI3VX0 $T=67200 194880 0 180 $X=65090 $Y=189760
X9622 1 2 211 1191 INJI3VX0 $T=71680 159040 1 180 $X=69570 $Y=158400
X9623 1 2 212 214 INJI3VX0 $T=70560 185920 1 0 $X=70130 $Y=180800
X9624 1 2 772 210 INJI3VX0 $T=75040 203840 0 180 $X=72930 $Y=198720
X9625 1 2 779 114 INJI3VX0 $T=83440 24640 0 0 $X=83010 $Y=24000
X9626 1 2 223 1419 INJI3VX0 $T=84000 33600 0 0 $X=83570 $Y=32960
X9627 1 2 762 1006 INJI3VX0 $T=94080 24640 1 180 $X=91970 $Y=24000
X9628 1 2 783 1418 INJI3VX0 $T=92960 42560 0 0 $X=92530 $Y=41920
X9629 1 2 241 786 INJI3VX0 $T=108640 33600 0 180 $X=106530 $Y=28480
X9630 1 2 245 793 INJI3VX0 $T=117040 24640 0 0 $X=116610 $Y=24000
X9631 1 2 801 1015 INJI3VX0 $T=123200 24640 0 0 $X=122770 $Y=24000
X9632 1 2 288 809 INJI3VX0 $T=136640 33600 0 0 $X=136210 $Y=32960
X9633 1 2 291 810 INJI3VX0 $T=139440 159040 0 0 $X=139010 $Y=158400
X9634 1 2 817 1420 INJI3VX0 $T=141680 24640 1 180 $X=139570 $Y=24000
X9635 1 2 1038 1342 INJI3VX0 $T=152880 123200 0 180 $X=150770 $Y=118080
X9636 1 2 1036 314 INJI3VX0 $T=154560 33600 1 180 $X=152450 $Y=32960
X9637 1 2 312 1221 INJI3VX0 $T=152880 123200 1 0 $X=152450 $Y=118080
X9638 1 2 367 1368 INJI3VX0 $T=164640 114240 1 180 $X=162530 $Y=113600
X9639 1 2 322 1421 INJI3VX0 $T=164640 24640 1 0 $X=164210 $Y=19520
X9640 1 2 334 341 INJI3VX0 $T=168000 24640 1 0 $X=167570 $Y=19520
X9641 1 2 348 324 INJI3VX0 $T=170800 123200 1 180 $X=168690 $Y=122560
X9642 1 2 382 310 INJI3VX0 $T=172480 176960 0 180 $X=170370 $Y=171840
X9643 1 2 304 351 INJI3VX0 $T=172480 114240 0 0 $X=172050 $Y=113600
X9644 1 2 358 313 INJI3VX0 $T=175840 176960 0 180 $X=173730 $Y=171840
X9645 1 2 355 842 INJI3VX0 $T=175840 203840 1 0 $X=175410 $Y=198720
X9646 1 2 360 1060 INJI3VX0 $T=178080 168000 0 0 $X=177650 $Y=167360
X9647 1 2 1055 369 INJI3VX0 $T=178640 194880 0 0 $X=178210 $Y=194240
X9648 1 2 121 1422 INJI3VX0 $T=183120 33600 1 0 $X=182690 $Y=28480
X9649 1 2 379 844 INJI3VX0 $T=183680 203840 0 0 $X=183250 $Y=203200
X9650 1 2 361 1431 INJI3VX0 $T=184240 176960 0 0 $X=183810 $Y=176320
X9651 1 2 847 1387 INJI3VX0 $T=190960 176960 0 0 $X=190530 $Y=176320
X9652 1 2 343 1238 INJI3VX0 $T=192080 185920 1 0 $X=191650 $Y=180800
X9653 1 2 852 1243 INJI3VX0 $T=204400 203840 0 180 $X=202290 $Y=198720
X9654 1 2 125 718 INJI3VX0 $T=203280 194880 0 0 $X=202850 $Y=194240
X9655 1 2 413 1077 INJI3VX0 $T=205520 33600 0 0 $X=205090 $Y=32960
X9656 1 2 398 412 INJI3VX0 $T=208880 42560 1 180 $X=206770 $Y=41920
X9657 1 2 319 1347 INJI3VX0 $T=208320 203840 0 0 $X=207890 $Y=203200
X9658 1 2 420 1079 INJI3VX0 $T=209440 176960 1 0 $X=209010 $Y=171840
X9659 1 2 416 1081 INJI3VX0 $T=209440 203840 1 0 $X=209010 $Y=198720
X9660 1 2 418 1434 INJI3VX0 $T=211120 159040 1 0 $X=210690 $Y=153920
X9661 1 2 549 1085 INJI3VX0 $T=215040 168000 1 0 $X=214610 $Y=162880
X9662 1 2 1080 132 INJI3VX0 $T=215600 185920 0 0 $X=215170 $Y=185280
X9663 1 2 453 856 INJI3VX0 $T=219520 185920 1 180 $X=217410 $Y=185280
X9664 1 2 428 1423 INJI3VX0 $T=219520 33600 1 0 $X=219090 $Y=28480
X9665 1 2 461 1330 INJI3VX0 $T=233520 33600 0 180 $X=231410 $Y=28480
X9666 1 2 1095 883 INJI3VX0 $T=241920 185920 0 0 $X=241490 $Y=185280
X9667 1 2 471 1424 INJI3VX0 $T=246960 24640 1 180 $X=244850 $Y=24000
X9668 1 2 888 448 INJI3VX0 $T=250320 185920 0 180 $X=248210 $Y=180800
X9669 1 2 456 472 INJI3VX0 $T=257040 185920 1 180 $X=254930 $Y=185280
X9670 1 2 470 1267 INJI3VX0 $T=257600 176960 1 0 $X=257170 $Y=171840
X9671 1 2 479 1111 INJI3VX0 $T=262640 194880 0 180 $X=260530 $Y=189760
X9672 1 2 485 1170 INJI3VX0 $T=264320 194880 0 180 $X=262210 $Y=189760
X9673 1 2 902 481 INJI3VX0 $T=265440 185920 0 180 $X=263330 $Y=180800
X9674 1 2 490 1112 INJI3VX0 $T=266000 194880 0 180 $X=263890 $Y=189760
X9675 1 2 100 492 INJI3VX0 $T=267680 194880 0 180 $X=265570 $Y=189760
X9676 1 2 497 1425 INJI3VX0 $T=269360 24640 1 180 $X=267250 $Y=24000
X9677 1 2 906 1256 INJI3VX0 $T=273280 194880 0 180 $X=271170 $Y=189760
X9678 1 2 501 1118 INJI3VX0 $T=272160 42560 0 0 $X=271730 $Y=41920
X9679 1 2 512 1426 INJI3VX0 $T=276640 33600 0 0 $X=276210 $Y=32960
X9680 1 2 903 523 INJI3VX0 $T=278880 185920 0 0 $X=278450 $Y=185280
X9681 1 2 920 1126 INJI3VX0 $T=295120 42560 0 0 $X=294690 $Y=41920
X9682 1 2 539 921 INJI3VX0 $T=297360 168000 1 0 $X=296930 $Y=162880
X9683 1 2 532 1427 INJI3VX0 $T=300720 24640 0 180 $X=298610 $Y=19520
X9684 1 2 137 567 INJI3VX0 $T=315280 33600 0 0 $X=314850 $Y=32960
X9685 1 2 1123 1132 INJI3VX0 $T=319760 159040 0 0 $X=319330 $Y=158400
X9686 1 2 589 931 INJI3VX0 $T=321440 168000 0 180 $X=319330 $Y=162880
X9687 1 2 1134 1133 INJI3VX0 $T=323680 24640 1 180 $X=321570 $Y=24000
X9688 1 2 594 937 INJI3VX0 $T=333760 33600 1 0 $X=333330 $Y=28480
X9689 1 2 139 612 INJI3VX0 $T=337680 176960 0 0 $X=337250 $Y=176320
X9690 1 2 140 1138 INJI3VX0 $T=340480 176960 1 0 $X=340050 $Y=171840
X9691 1 2 1145 947 INJI3VX0 $T=344400 185920 0 0 $X=343970 $Y=185280
X9692 1 2 587 948 INJI3VX0 $T=345520 194880 1 0 $X=345090 $Y=189760
X9693 1 2 623 618 INJI3VX0 $T=347760 168000 0 180 $X=345650 $Y=162880
X9694 1 2 1149 624 INJI3VX0 $T=346640 51520 1 0 $X=346210 $Y=46400
X9695 1 2 630 627 INJI3VX0 $T=347760 176960 1 0 $X=347330 $Y=171840
X9696 1 2 622 619 INJI3VX0 $T=348320 212800 1 0 $X=347890 $Y=207680
X9697 1 2 636 104 INJI3VX0 $T=362880 176960 0 180 $X=360770 $Y=171840
X9698 1 2 954 1146 INJI3VX0 $T=364560 176960 1 180 $X=362450 $Y=176320
X9699 1 2 143 1428 INJI3VX0 $T=367920 33600 1 180 $X=365810 $Y=32960
X9700 1 2 647 648 INJI3VX0 $T=374640 24640 0 0 $X=374210 $Y=24000
X9701 1 2 650 1309 INJI3VX0 $T=375200 42560 1 0 $X=374770 $Y=37440
X9702 1 2 661 667 INJI3VX0 $T=381360 141120 0 180 $X=379250 $Y=136000
X9703 1 2 670 664 INJI3VX0 $T=384160 123200 1 180 $X=382050 $Y=122560
X9704 1 2 659 673 INJI3VX0 $T=385840 132160 0 0 $X=385410 $Y=131520
X9705 1 2 693 1312 INJI3VX0 $T=389200 123200 1 0 $X=388770 $Y=118080
X9706 1 2 1159 679 INJI3VX0 $T=390880 150080 1 180 $X=388770 $Y=149440
X9707 1 2 687 1166 INJI3VX0 $T=392560 123200 0 0 $X=392130 $Y=122560
X9708 1 2 1165 685 INJI3VX0 $T=394240 159040 1 180 $X=392130 $Y=158400
X9709 1 2 694 1429 INJI3VX0 $T=397040 24640 1 180 $X=394930 $Y=24000
X9710 1 2 683 966 INJI3VX0 $T=395920 159040 1 0 $X=395490 $Y=153920
X9711 1 2 1413 688 INJI3VX0 $T=398160 141120 0 180 $X=396050 $Y=136000
X9712 1 2 971 684 INJI3VX0 $T=405440 33600 1 180 $X=403330 $Y=32960
X9713 1 2 761 1370 750 195 NO3I1JI3VX1 $T=57120 168000 1 0 $X=56690 $Y=162880
X9714 1 2 840 1412 122 1067 NO3I1JI3VX1 $T=187040 185920 1 0 $X=186610 $Y=180800
X9715 1 2 1246 286 304 1433 NO3I1JI3VX1 $T=206080 159040 0 180 $X=201170 $Y=153920
X9716 1 2 1105 869 469 1432 NO3I1JI3VX1 $T=254240 168000 1 0 $X=253810 $Y=162880
X9717 1 2 575 1396 928 564 NO3I1JI3VX1 $T=319760 168000 0 180 $X=314850 $Y=162880
X9718 1 2 DECAP25JI3V $T=20160 24640 1 0 $X=19730 $Y=19520
X9719 1 2 DECAP25JI3V $T=20160 24640 0 0 $X=19730 $Y=24000
X9720 1 2 DECAP25JI3V $T=20160 33600 1 0 $X=19730 $Y=28480
X9721 1 2 DECAP25JI3V $T=20160 42560 1 0 $X=19730 $Y=37440
X9722 1 2 DECAP25JI3V $T=20160 42560 0 0 $X=19730 $Y=41920
X9723 1 2 DECAP25JI3V $T=20160 51520 1 0 $X=19730 $Y=46400
X9724 1 2 DECAP25JI3V $T=20160 51520 0 0 $X=19730 $Y=50880
X9725 1 2 DECAP25JI3V $T=20160 60480 1 0 $X=19730 $Y=55360
X9726 1 2 DECAP25JI3V $T=20160 60480 0 0 $X=19730 $Y=59840
X9727 1 2 DECAP25JI3V $T=20160 69440 1 0 $X=19730 $Y=64320
X9728 1 2 DECAP25JI3V $T=20160 69440 0 0 $X=19730 $Y=68800
X9729 1 2 DECAP25JI3V $T=20160 78400 1 0 $X=19730 $Y=73280
X9730 1 2 DECAP25JI3V $T=20160 78400 0 0 $X=19730 $Y=77760
X9731 1 2 DECAP25JI3V $T=20160 87360 1 0 $X=19730 $Y=82240
X9732 1 2 DECAP25JI3V $T=20160 87360 0 0 $X=19730 $Y=86720
X9733 1 2 DECAP25JI3V $T=20160 96320 1 0 $X=19730 $Y=91200
X9734 1 2 DECAP25JI3V $T=20160 141120 0 0 $X=19730 $Y=140480
X9735 1 2 DECAP25JI3V $T=20160 194880 0 0 $X=19730 $Y=194240
X9736 1 2 DECAP25JI3V $T=20160 203840 1 0 $X=19730 $Y=198720
X9737 1 2 DECAP25JI3V $T=20160 203840 0 0 $X=19730 $Y=203200
X9738 1 2 DECAP25JI3V $T=20160 212800 1 0 $X=19730 $Y=207680
X9739 1 2 DECAP25JI3V $T=20160 212800 0 0 $X=19730 $Y=212160
X9740 1 2 DECAP25JI3V $T=34160 33600 1 0 $X=33730 $Y=28480
X9741 1 2 DECAP25JI3V $T=34160 60480 0 0 $X=33730 $Y=59840
X9742 1 2 DECAP25JI3V $T=34160 87360 0 0 $X=33730 $Y=86720
X9743 1 2 DECAP25JI3V $T=34160 203840 1 0 $X=33730 $Y=198720
X9744 1 2 DECAP25JI3V $T=34160 212800 1 0 $X=33730 $Y=207680
X9745 1 2 DECAP25JI3V $T=34160 212800 0 0 $X=33730 $Y=212160
X9746 1 2 DECAP25JI3V $T=48160 87360 0 0 $X=47730 $Y=86720
X9747 1 2 DECAP25JI3V $T=48160 212800 0 0 $X=47730 $Y=212160
X9748 1 2 DECAP25JI3V $T=57120 132160 0 0 $X=56690 $Y=131520
X9749 1 2 DECAP25JI3V $T=80080 123200 1 0 $X=79650 $Y=118080
X9750 1 2 DECAP25JI3V $T=85680 96320 0 0 $X=85250 $Y=95680
X9751 1 2 DECAP25JI3V $T=86240 87360 0 0 $X=85810 $Y=86720
X9752 1 2 DECAP25JI3V $T=86240 105280 1 0 $X=85810 $Y=100160
X9753 1 2 DECAP25JI3V $T=89040 114240 0 0 $X=88610 $Y=113600
X9754 1 2 DECAP25JI3V $T=93520 105280 0 0 $X=93090 $Y=104640
X9755 1 2 DECAP25JI3V $T=110880 87360 0 180 $X=96450 $Y=82240
X9756 1 2 DECAP25JI3V $T=215040 114240 0 0 $X=214610 $Y=113600
X9757 1 2 DECAP25JI3V $T=223440 123200 0 0 $X=223010 $Y=122560
X9758 1 2 DECAP25JI3V $T=231840 96320 1 0 $X=231410 $Y=91200
X9759 1 2 DECAP25JI3V $T=257600 114240 0 0 $X=257170 $Y=113600
X9760 1 2 DECAP25JI3V $T=271600 114240 0 0 $X=271170 $Y=113600
X9761 1 2 DECAP25JI3V $T=295120 78400 0 0 $X=294690 $Y=77760
X9762 1 2 DECAP25JI3V $T=308000 132160 0 0 $X=307570 $Y=131520
X9763 1 2 DECAP25JI3V $T=312480 105280 0 0 $X=312050 $Y=104640
X9764 1 2 DECAP25JI3V $T=313040 194880 0 0 $X=312610 $Y=194240
X9765 1 2 DECAP25JI3V $T=318080 123200 0 0 $X=317650 $Y=122560
X9766 1 2 DECAP25JI3V $T=333760 114240 1 0 $X=333330 $Y=109120
X9767 1 2 DECAP25JI3V $T=336000 105280 1 0 $X=335570 $Y=100160
X9768 1 2 DECAP25JI3V $T=338240 87360 1 0 $X=337810 $Y=82240
X9769 1 2 DECAP25JI3V $T=350000 212800 1 0 $X=349570 $Y=207680
X9770 1 2 DECAP25JI3V $T=351120 203840 0 0 $X=350690 $Y=203200
X9771 1 2 DECAP25JI3V $T=352240 212800 0 0 $X=351810 $Y=212160
X9772 1 2 DECAP25JI3V $T=352800 203840 1 0 $X=352370 $Y=198720
X9773 1 2 DECAP25JI3V $T=364000 212800 1 0 $X=363570 $Y=207680
X9774 1 2 DECAP25JI3V $T=365120 203840 0 0 $X=364690 $Y=203200
X9775 1 2 DECAP25JI3V $T=366240 212800 0 0 $X=365810 $Y=212160
X9776 1 2 DECAP25JI3V $T=366800 203840 1 0 $X=366370 $Y=198720
X9777 1 2 DECAP25JI3V $T=370160 194880 1 0 $X=369730 $Y=189760
X9778 1 2 DECAP25JI3V $T=371280 194880 0 0 $X=370850 $Y=194240
X9779 1 2 DECAP25JI3V $T=378000 212800 1 0 $X=377570 $Y=207680
X9780 1 2 DECAP25JI3V $T=379120 185920 0 0 $X=378690 $Y=185280
X9781 1 2 DECAP25JI3V $T=379120 203840 0 0 $X=378690 $Y=203200
X9782 1 2 DECAP25JI3V $T=380240 212800 0 0 $X=379810 $Y=212160
X9783 1 2 DECAP25JI3V $T=380800 176960 0 0 $X=380370 $Y=176320
X9784 1 2 DECAP25JI3V $T=380800 203840 1 0 $X=380370 $Y=198720
X9785 1 2 DECAP25JI3V $T=381360 176960 1 0 $X=380930 $Y=171840
X9786 1 2 DECAP25JI3V $T=384160 194880 1 0 $X=383730 $Y=189760
X9787 1 2 DECAP25JI3V $T=385280 194880 0 0 $X=384850 $Y=194240
X9788 1 2 DECAP25JI3V $T=389200 185920 1 0 $X=388770 $Y=180800
X9789 1 2 DECAP25JI3V $T=392000 212800 1 0 $X=391570 $Y=207680
X9790 1 2 DECAP25JI3V $T=393120 185920 0 0 $X=392690 $Y=185280
X9791 1 2 DECAP25JI3V $T=393120 203840 0 0 $X=392690 $Y=203200
X9792 1 2 DECAP25JI3V $T=394240 212800 0 0 $X=393810 $Y=212160
X9793 1 2 DECAP25JI3V $T=394800 176960 0 0 $X=394370 $Y=176320
X9794 1 2 DECAP25JI3V $T=394800 203840 1 0 $X=394370 $Y=198720
X9795 1 2 DECAP25JI3V $T=395360 176960 1 0 $X=394930 $Y=171840
X9796 1 2 DECAP25JI3V $T=398160 194880 1 0 $X=397730 $Y=189760
X9797 1 2 DECAP25JI3V $T=398720 141120 0 0 $X=398290 $Y=140480
X9798 1 2 DECAP25JI3V $T=398720 150080 1 0 $X=398290 $Y=144960
X9799 1 2 DECAP25JI3V $T=399280 194880 0 0 $X=398850 $Y=194240
X9800 1 2 DECAP25JI3V $T=399840 159040 0 0 $X=399410 $Y=158400
X9801 1 2 DECAP25JI3V $T=400400 78400 0 0 $X=399970 $Y=77760
X9802 1 2 DECAP25JI3V $T=400400 96320 0 0 $X=399970 $Y=95680
X9803 1 2 DECAP25JI3V $T=414400 168000 0 180 $X=399970 $Y=162880
X9804 1 2 DECAP25JI3V $T=402080 141120 1 0 $X=401650 $Y=136000
X9805 1 2 DECAP25JI3V $T=403200 185920 1 0 $X=402770 $Y=180800
X9806 1 2 DECAP25JI3V $T=404320 159040 1 0 $X=403890 $Y=153920
X9807 1 2 DECAP25JI3V $T=406000 24640 1 0 $X=405570 $Y=19520
X9808 1 2 DECAP25JI3V $T=406000 212800 1 0 $X=405570 $Y=207680
X9809 1 2 DECAP25JI3V $T=406560 105280 0 0 $X=406130 $Y=104640
X9810 1 2 DECAP25JI3V $T=406560 114240 1 0 $X=406130 $Y=109120
X9811 1 2 DECAP25JI3V $T=407120 185920 0 0 $X=406690 $Y=185280
X9812 1 2 DECAP25JI3V $T=407120 203840 0 0 $X=406690 $Y=203200
X9813 1 2 DECAP25JI3V $T=407680 168000 0 0 $X=407250 $Y=167360
X9814 1 2 DECAP25JI3V $T=408800 150080 0 0 $X=408370 $Y=149440
X9815 1 2 DECAP25JI3V $T=408800 176960 0 0 $X=408370 $Y=176320
X9816 1 2 DECAP25JI3V $T=408800 203840 1 0 $X=408370 $Y=198720
X9817 1 2 DECAP25JI3V $T=409360 24640 0 0 $X=408930 $Y=24000
X9818 1 2 DECAP25JI3V $T=409360 176960 1 0 $X=408930 $Y=171840
X9819 1 2 DECAP25JI3V $T=409920 132160 1 0 $X=409490 $Y=127040
X9820 1 2 DECAP25JI3V $T=412720 132160 0 0 $X=412290 $Y=131520
X9821 1 2 DECAP25JI3V $T=412720 141120 0 0 $X=412290 $Y=140480
X9822 1 2 DECAP25JI3V $T=412720 150080 1 0 $X=412290 $Y=144960
X9823 1 2 DECAP25JI3V $T=413280 42560 1 0 $X=412850 $Y=37440
X9824 1 2 DECAP25JI3V $T=413280 60480 0 0 $X=412850 $Y=59840
X9825 1 2 DECAP25JI3V $T=413280 69440 1 0 $X=412850 $Y=64320
X9826 1 2 DECAP25JI3V $T=413280 69440 0 0 $X=412850 $Y=68800
X9827 1 2 DECAP25JI3V $T=413280 105280 1 0 $X=412850 $Y=100160
X9828 1 2 DECAP25JI3V $T=413280 194880 0 0 $X=412850 $Y=194240
X9829 1 2 DECAP25JI3V $T=414400 78400 0 0 $X=413970 $Y=77760
X9830 1 2 DECAP25JI3V $T=414400 96320 0 0 $X=413970 $Y=95680
X9831 1 2 DECAP25JI3V $T=414400 168000 1 0 $X=413970 $Y=162880
X9832 1 2 DECAP25JI3V $T=417200 185920 1 0 $X=416770 $Y=180800
X9833 1 2 DECAP25JI3V $T=418320 159040 1 0 $X=417890 $Y=153920
X9834 1 2 DECAP25JI3V $T=421120 185920 0 0 $X=420690 $Y=185280
X9835 1 2 DECAP25JI3V $T=421120 203840 0 0 $X=420690 $Y=203200
X9836 1 2 DECAP15JI3V $T=20160 33600 0 0 $X=19730 $Y=32960
X9837 1 2 DECAP15JI3V $T=20160 96320 0 0 $X=19730 $Y=95680
X9838 1 2 DECAP15JI3V $T=20160 141120 1 0 $X=19730 $Y=136000
X9839 1 2 DECAP15JI3V $T=34160 24640 1 0 $X=33730 $Y=19520
X9840 1 2 DECAP15JI3V $T=34160 60480 1 0 $X=33730 $Y=55360
X9841 1 2 DECAP15JI3V $T=34160 69440 0 0 $X=33730 $Y=68800
X9842 1 2 DECAP15JI3V $T=34160 78400 1 0 $X=33730 $Y=73280
X9843 1 2 DECAP15JI3V $T=34160 203840 0 0 $X=33730 $Y=203200
X9844 1 2 DECAP15JI3V $T=48160 60480 0 0 $X=47730 $Y=59840
X9845 1 2 DECAP15JI3V $T=48160 212800 1 0 $X=47730 $Y=207680
X9846 1 2 DECAP15JI3V $T=54880 114240 0 0 $X=54450 $Y=113600
X9847 1 2 DECAP15JI3V $T=61040 69440 1 0 $X=60610 $Y=64320
X9848 1 2 DECAP15JI3V $T=62720 69440 0 0 $X=62290 $Y=68800
X9849 1 2 DECAP15JI3V $T=62720 78400 1 0 $X=62290 $Y=73280
X9850 1 2 DECAP15JI3V $T=80080 132160 1 0 $X=79650 $Y=127040
X9851 1 2 DECAP15JI3V $T=84000 123200 0 0 $X=83570 $Y=122560
X9852 1 2 DECAP15JI3V $T=86800 96320 1 0 $X=86370 $Y=91200
X9853 1 2 DECAP15JI3V $T=90160 185920 1 0 $X=89730 $Y=180800
X9854 1 2 DECAP15JI3V $T=90160 212800 1 0 $X=89730 $Y=207680
X9855 1 2 DECAP15JI3V $T=91280 150080 0 0 $X=90850 $Y=149440
X9856 1 2 DECAP15JI3V $T=91840 159040 1 0 $X=91410 $Y=153920
X9857 1 2 DECAP15JI3V $T=94080 123200 1 0 $X=93650 $Y=118080
X9858 1 2 DECAP15JI3V $T=95200 69440 0 0 $X=94770 $Y=68800
X9859 1 2 DECAP15JI3V $T=99680 96320 0 0 $X=99250 $Y=95680
X9860 1 2 DECAP15JI3V $T=100240 78400 0 0 $X=99810 $Y=77760
X9861 1 2 DECAP15JI3V $T=103040 114240 0 0 $X=102610 $Y=113600
X9862 1 2 DECAP15JI3V $T=108080 96320 0 0 $X=107650 $Y=95680
X9863 1 2 DECAP15JI3V $T=123200 78400 1 0 $X=122770 $Y=73280
X9864 1 2 DECAP15JI3V $T=128240 194880 1 0 $X=127810 $Y=189760
X9865 1 2 DECAP15JI3V $T=137760 159040 1 180 $X=128930 $Y=158400
X9866 1 2 DECAP15JI3V $T=131600 78400 0 0 $X=131170 $Y=77760
X9867 1 2 DECAP15JI3V $T=151200 168000 1 0 $X=150770 $Y=162880
X9868 1 2 DECAP15JI3V $T=162960 78400 0 0 $X=162530 $Y=77760
X9869 1 2 DECAP15JI3V $T=210000 87360 1 0 $X=209570 $Y=82240
X9870 1 2 DECAP15JI3V $T=215600 42560 0 0 $X=215170 $Y=41920
X9871 1 2 DECAP15JI3V $T=215600 51520 1 0 $X=215170 $Y=46400
X9872 1 2 DECAP15JI3V $T=223440 33600 0 0 $X=223010 $Y=32960
X9873 1 2 DECAP15JI3V $T=223440 69440 0 0 $X=223010 $Y=68800
X9874 1 2 DECAP15JI3V $T=223440 78400 1 0 $X=223010 $Y=73280
X9875 1 2 DECAP15JI3V $T=223440 96320 1 0 $X=223010 $Y=91200
X9876 1 2 DECAP15JI3V $T=223440 105280 1 0 $X=223010 $Y=100160
X9877 1 2 DECAP15JI3V $T=223440 114240 1 0 $X=223010 $Y=109120
X9878 1 2 DECAP15JI3V $T=229040 114240 0 0 $X=228610 $Y=113600
X9879 1 2 DECAP15JI3V $T=258720 78400 0 0 $X=258290 $Y=77760
X9880 1 2 DECAP15JI3V $T=267120 212800 1 0 $X=266690 $Y=207680
X9881 1 2 DECAP15JI3V $T=268800 212800 0 0 $X=268370 $Y=212160
X9882 1 2 DECAP15JI3V $T=276640 105280 1 0 $X=276210 $Y=100160
X9883 1 2 DECAP15JI3V $T=279440 42560 0 0 $X=279010 $Y=41920
X9884 1 2 DECAP15JI3V $T=280560 185920 0 0 $X=280130 $Y=185280
X9885 1 2 DECAP15JI3V $T=294560 96320 0 0 $X=294130 $Y=95680
X9886 1 2 DECAP15JI3V $T=298480 194880 1 0 $X=298050 $Y=189760
X9887 1 2 DECAP15JI3V $T=300720 114240 1 0 $X=300290 $Y=109120
X9888 1 2 DECAP15JI3V $T=327600 203840 0 0 $X=327170 $Y=203200
X9889 1 2 DECAP15JI3V $T=336000 96320 0 0 $X=335570 $Y=95680
X9890 1 2 DECAP15JI3V $T=337120 96320 1 0 $X=336690 $Y=91200
X9891 1 2 DECAP15JI3V $T=337120 114240 0 0 $X=336690 $Y=113600
X9892 1 2 DECAP15JI3V $T=344960 194880 0 0 $X=344530 $Y=194240
X9893 1 2 DECAP15JI3V $T=350000 105280 1 0 $X=349570 $Y=100160
X9894 1 2 DECAP15JI3V $T=350000 185920 1 0 $X=349570 $Y=180800
X9895 1 2 DECAP15JI3V $T=351680 51520 1 0 $X=351250 $Y=46400
X9896 1 2 DECAP15JI3V $T=351680 69440 0 0 $X=351250 $Y=68800
X9897 1 2 DECAP15JI3V $T=351680 78400 1 0 $X=351250 $Y=73280
X9898 1 2 DECAP15JI3V $T=352240 24640 0 0 $X=351810 $Y=24000
X9899 1 2 DECAP15JI3V $T=381920 141120 1 180 $X=373090 $Y=140480
X9900 1 2 DECAP15JI3V $T=388640 96320 0 180 $X=379810 $Y=91200
X9901 1 2 DECAP15JI3V $T=380800 185920 1 0 $X=380370 $Y=180800
X9902 1 2 DECAP15JI3V $T=381360 78400 1 0 $X=380930 $Y=73280
X9903 1 2 DECAP15JI3V $T=416640 33600 0 180 $X=407810 $Y=28480
X9904 1 2 DECAP15JI3V $T=408240 212800 0 0 $X=407810 $Y=212160
X9905 1 2 DECAP15JI3V $T=411040 114240 0 0 $X=410610 $Y=113600
X9906 1 2 DECAP15JI3V $T=412160 194880 1 0 $X=411730 $Y=189760
X9907 1 2 DECAP15JI3V $T=413280 33600 0 0 $X=412850 $Y=32960
X9908 1 2 DECAP15JI3V $T=413280 60480 1 0 $X=412850 $Y=55360
X9909 1 2 DECAP15JI3V $T=416080 123200 1 0 $X=415650 $Y=118080
X9910 1 2 DECAP15JI3V $T=416080 141120 1 0 $X=415650 $Y=136000
X9911 1 2 DECAP15JI3V $T=418880 42560 0 0 $X=418450 $Y=41920
X9912 1 2 DECAP15JI3V $T=418880 51520 1 0 $X=418450 $Y=46400
X9913 1 2 DECAP15JI3V $T=418880 51520 0 0 $X=418450 $Y=50880
X9914 1 2 DECAP15JI3V $T=420000 24640 1 0 $X=419570 $Y=19520
X9915 1 2 DECAP15JI3V $T=420000 212800 1 0 $X=419570 $Y=207680
X9916 1 2 DECAP15JI3V $T=422800 150080 0 0 $X=422370 $Y=149440
X9917 1 2 DECAP15JI3V $T=422800 176960 0 0 $X=422370 $Y=176320
X9918 1 2 DECAP15JI3V $T=422800 203840 1 0 $X=422370 $Y=198720
X9919 1 2 DECAP15JI3V $T=423920 132160 1 0 $X=423490 $Y=127040
X9920 1 2 DECAP15JI3V $T=426720 132160 0 0 $X=426290 $Y=131520
X9921 1 2 DECAP15JI3V $T=426720 141120 0 0 $X=426290 $Y=140480
X9922 1 2 DECAP15JI3V $T=426720 150080 1 0 $X=426290 $Y=144960
X9923 1 2 DECAP7JI3V $T=20160 105280 1 0 $X=19730 $Y=100160
X9924 1 2 DECAP7JI3V $T=20160 150080 0 0 $X=19730 $Y=149440
X9925 1 2 DECAP7JI3V $T=20160 168000 1 0 $X=19730 $Y=162880
X9926 1 2 DECAP7JI3V $T=20160 168000 0 0 $X=19730 $Y=167360
X9927 1 2 DECAP7JI3V $T=25760 114240 0 0 $X=25330 $Y=113600
X9928 1 2 DECAP7JI3V $T=25760 123200 1 0 $X=25330 $Y=118080
X9929 1 2 DECAP7JI3V $T=25760 176960 0 0 $X=25330 $Y=176320
X9930 1 2 DECAP7JI3V $T=28560 33600 0 0 $X=28130 $Y=32960
X9931 1 2 DECAP7JI3V $T=28560 96320 0 0 $X=28130 $Y=95680
X9932 1 2 DECAP7JI3V $T=32480 33600 0 0 $X=32050 $Y=32960
X9933 1 2 DECAP7JI3V $T=34160 42560 1 0 $X=33730 $Y=37440
X9934 1 2 DECAP7JI3V $T=34160 42560 0 0 $X=33730 $Y=41920
X9935 1 2 DECAP7JI3V $T=34160 51520 1 0 $X=33730 $Y=46400
X9936 1 2 DECAP7JI3V $T=34160 51520 0 0 $X=33730 $Y=50880
X9937 1 2 DECAP7JI3V $T=34160 69440 1 0 $X=33730 $Y=64320
X9938 1 2 DECAP7JI3V $T=34160 78400 0 0 $X=33730 $Y=77760
X9939 1 2 DECAP7JI3V $T=34160 96320 1 0 $X=33730 $Y=91200
X9940 1 2 DECAP7JI3V $T=36400 33600 0 0 $X=35970 $Y=32960
X9941 1 2 DECAP7JI3V $T=36960 123200 1 0 $X=36530 $Y=118080
X9942 1 2 DECAP7JI3V $T=38080 42560 1 0 $X=37650 $Y=37440
X9943 1 2 DECAP7JI3V $T=38080 42560 0 0 $X=37650 $Y=41920
X9944 1 2 DECAP7JI3V $T=38080 51520 1 0 $X=37650 $Y=46400
X9945 1 2 DECAP7JI3V $T=38080 51520 0 0 $X=37650 $Y=50880
X9946 1 2 DECAP7JI3V $T=38080 69440 1 0 $X=37650 $Y=64320
X9947 1 2 DECAP7JI3V $T=38080 96320 1 0 $X=37650 $Y=91200
X9948 1 2 DECAP7JI3V $T=39760 24640 0 0 $X=39330 $Y=24000
X9949 1 2 DECAP7JI3V $T=39760 194880 0 0 $X=39330 $Y=194240
X9950 1 2 DECAP7JI3V $T=40320 33600 0 0 $X=39890 $Y=32960
X9951 1 2 DECAP7JI3V $T=42000 69440 1 0 $X=41570 $Y=64320
X9952 1 2 DECAP7JI3V $T=42560 24640 1 0 $X=42130 $Y=19520
X9953 1 2 DECAP7JI3V $T=42560 203840 0 0 $X=42130 $Y=203200
X9954 1 2 DECAP7JI3V $T=43680 24640 0 0 $X=43250 $Y=24000
X9955 1 2 DECAP7JI3V $T=43680 194880 0 0 $X=43250 $Y=194240
X9956 1 2 DECAP7JI3V $T=46480 24640 1 0 $X=46050 $Y=19520
X9957 1 2 DECAP7JI3V $T=46480 203840 0 0 $X=46050 $Y=203200
X9958 1 2 DECAP7JI3V $T=47600 24640 0 0 $X=47170 $Y=24000
X9959 1 2 DECAP7JI3V $T=50400 24640 1 0 $X=49970 $Y=19520
X9960 1 2 DECAP7JI3V $T=50400 203840 0 0 $X=49970 $Y=203200
X9961 1 2 DECAP7JI3V $T=51520 24640 0 0 $X=51090 $Y=24000
X9962 1 2 DECAP7JI3V $T=54320 203840 0 0 $X=53890 $Y=203200
X9963 1 2 DECAP7JI3V $T=56560 60480 0 0 $X=56130 $Y=59840
X9964 1 2 DECAP7JI3V $T=56560 212800 1 0 $X=56130 $Y=207680
X9965 1 2 DECAP7JI3V $T=59920 51520 0 0 $X=59490 $Y=50880
X9966 1 2 DECAP7JI3V $T=60480 212800 1 0 $X=60050 $Y=207680
X9967 1 2 DECAP7JI3V $T=62160 212800 0 0 $X=61730 $Y=212160
X9968 1 2 DECAP7JI3V $T=62720 194880 0 0 $X=62290 $Y=194240
X9969 1 2 DECAP7JI3V $T=63280 114240 1 0 $X=62850 $Y=109120
X9970 1 2 DECAP7JI3V $T=64400 212800 1 0 $X=63970 $Y=207680
X9971 1 2 DECAP7JI3V $T=66080 212800 0 0 $X=65650 $Y=212160
X9972 1 2 DECAP7JI3V $T=67200 114240 1 0 $X=66770 $Y=109120
X9973 1 2 DECAP7JI3V $T=68320 212800 1 0 $X=67890 $Y=207680
X9974 1 2 DECAP7JI3V $T=70000 212800 0 0 $X=69570 $Y=212160
X9975 1 2 DECAP7JI3V $T=71120 78400 1 0 $X=70690 $Y=73280
X9976 1 2 DECAP7JI3V $T=71120 114240 1 0 $X=70690 $Y=109120
X9977 1 2 DECAP7JI3V $T=71120 132160 0 0 $X=70690 $Y=131520
X9978 1 2 DECAP7JI3V $T=80640 185920 0 0 $X=80210 $Y=185280
X9979 1 2 DECAP7JI3V $T=88480 132160 1 0 $X=88050 $Y=127040
X9980 1 2 DECAP7JI3V $T=90720 194880 0 0 $X=90290 $Y=194240
X9981 1 2 DECAP7JI3V $T=91280 185920 0 0 $X=90850 $Y=185280
X9982 1 2 DECAP7JI3V $T=92400 123200 0 0 $X=91970 $Y=122560
X9983 1 2 DECAP7JI3V $T=92400 132160 1 0 $X=91970 $Y=127040
X9984 1 2 DECAP7JI3V $T=93520 60480 0 0 $X=93090 $Y=59840
X9985 1 2 DECAP7JI3V $T=94640 42560 1 0 $X=94210 $Y=37440
X9986 1 2 DECAP7JI3V $T=94640 42560 0 0 $X=94210 $Y=41920
X9987 1 2 DECAP7JI3V $T=94640 194880 0 0 $X=94210 $Y=194240
X9988 1 2 DECAP7JI3V $T=95200 33600 1 0 $X=94770 $Y=28480
X9989 1 2 DECAP7JI3V $T=95200 69440 1 0 $X=94770 $Y=64320
X9990 1 2 DECAP7JI3V $T=95200 78400 1 0 $X=94770 $Y=73280
X9991 1 2 DECAP7JI3V $T=95200 96320 1 0 $X=94770 $Y=91200
X9992 1 2 DECAP7JI3V $T=95200 114240 1 0 $X=94770 $Y=109120
X9993 1 2 DECAP7JI3V $T=95200 132160 0 0 $X=94770 $Y=131520
X9994 1 2 DECAP7JI3V $T=95200 185920 0 0 $X=94770 $Y=185280
X9995 1 2 DECAP7JI3V $T=95200 203840 0 0 $X=94770 $Y=203200
X9996 1 2 DECAP7JI3V $T=96320 123200 0 0 $X=95890 $Y=122560
X9997 1 2 DECAP7JI3V $T=96320 132160 1 0 $X=95890 $Y=127040
X9998 1 2 DECAP7JI3V $T=96320 176960 1 0 $X=95890 $Y=171840
X9999 1 2 DECAP7JI3V $T=99120 33600 1 0 $X=98690 $Y=28480
X10000 1 2 DECAP7JI3V $T=99120 69440 1 0 $X=98690 $Y=64320
X10001 1 2 DECAP7JI3V $T=99120 78400 1 0 $X=98690 $Y=73280
X10002 1 2 DECAP7JI3V $T=99120 96320 1 0 $X=98690 $Y=91200
X10003 1 2 DECAP7JI3V $T=99120 114240 1 0 $X=98690 $Y=109120
X10004 1 2 DECAP7JI3V $T=99120 132160 0 0 $X=98690 $Y=131520
X10005 1 2 DECAP7JI3V $T=99120 185920 0 0 $X=98690 $Y=185280
X10006 1 2 DECAP7JI3V $T=99120 203840 0 0 $X=98690 $Y=203200
X10007 1 2 DECAP7JI3V $T=99680 150080 0 0 $X=99250 $Y=149440
X10008 1 2 DECAP7JI3V $T=100240 87360 0 0 $X=99810 $Y=86720
X10009 1 2 DECAP7JI3V $T=100240 176960 1 0 $X=99810 $Y=171840
X10010 1 2 DECAP7JI3V $T=100800 159040 0 0 $X=100370 $Y=158400
X10011 1 2 DECAP7JI3V $T=103040 33600 1 0 $X=102610 $Y=28480
X10012 1 2 DECAP7JI3V $T=103040 96320 1 0 $X=102610 $Y=91200
X10013 1 2 DECAP7JI3V $T=103040 114240 1 0 $X=102610 $Y=109120
X10014 1 2 DECAP7JI3V $T=104160 87360 0 0 $X=103730 $Y=86720
X10015 1 2 DECAP7JI3V $T=104720 159040 0 0 $X=104290 $Y=158400
X10016 1 2 DECAP7JI3V $T=105840 194880 1 0 $X=105410 $Y=189760
X10017 1 2 DECAP7JI3V $T=106960 96320 1 0 $X=106530 $Y=91200
X10018 1 2 DECAP7JI3V $T=106960 114240 1 0 $X=106530 $Y=109120
X10019 1 2 DECAP7JI3V $T=111440 114240 0 0 $X=111010 $Y=113600
X10020 1 2 DECAP7JI3V $T=116480 96320 0 0 $X=116050 $Y=95680
X10021 1 2 DECAP7JI3V $T=123200 69440 1 0 $X=122770 $Y=64320
X10022 1 2 DECAP7JI3V $T=128240 105280 0 180 $X=123890 $Y=100160
X10023 1 2 DECAP7JI3V $T=127120 69440 1 0 $X=126690 $Y=64320
X10024 1 2 DECAP7JI3V $T=132160 69440 0 0 $X=131730 $Y=68800
X10025 1 2 DECAP7JI3V $T=132160 87360 0 0 $X=131730 $Y=86720
X10026 1 2 DECAP7JI3V $T=135520 212800 0 0 $X=135090 $Y=212160
X10027 1 2 DECAP7JI3V $T=136080 87360 0 0 $X=135650 $Y=86720
X10028 1 2 DECAP7JI3V $T=138320 33600 0 0 $X=137890 $Y=32960
X10029 1 2 DECAP7JI3V $T=151760 78400 1 0 $X=151330 $Y=73280
X10030 1 2 DECAP7JI3V $T=155680 78400 1 0 $X=155250 $Y=73280
X10031 1 2 DECAP7JI3V $T=155680 203840 1 0 $X=155250 $Y=198720
X10032 1 2 DECAP7JI3V $T=158480 87360 1 0 $X=158050 $Y=82240
X10033 1 2 DECAP7JI3V $T=159600 168000 1 0 $X=159170 $Y=162880
X10034 1 2 DECAP7JI3V $T=162400 33600 0 0 $X=161970 $Y=32960
X10035 1 2 DECAP7JI3V $T=162960 60480 0 0 $X=162530 $Y=59840
X10036 1 2 DECAP7JI3V $T=166320 168000 0 0 $X=165890 $Y=167360
X10037 1 2 DECAP7JI3V $T=166880 60480 0 0 $X=166450 $Y=59840
X10038 1 2 DECAP7JI3V $T=169680 24640 1 0 $X=169250 $Y=19520
X10039 1 2 DECAP7JI3V $T=170240 168000 0 0 $X=169810 $Y=167360
X10040 1 2 DECAP7JI3V $T=170800 60480 0 0 $X=170370 $Y=59840
X10041 1 2 DECAP7JI3V $T=171360 78400 0 0 $X=170930 $Y=77760
X10042 1 2 DECAP7JI3V $T=178080 168000 1 180 $X=173730 $Y=167360
X10043 1 2 DECAP7JI3V $T=174720 60480 0 0 $X=174290 $Y=59840
X10044 1 2 DECAP7JI3V $T=175280 78400 0 0 $X=174850 $Y=77760
X10045 1 2 DECAP7JI3V $T=179200 78400 0 0 $X=178770 $Y=77760
X10046 1 2 DECAP7JI3V $T=184240 69440 0 0 $X=183810 $Y=68800
X10047 1 2 DECAP7JI3V $T=184800 194880 1 0 $X=184370 $Y=189760
X10048 1 2 DECAP7JI3V $T=197680 33600 0 0 $X=197250 $Y=32960
X10049 1 2 DECAP7JI3V $T=197680 60480 1 0 $X=197250 $Y=55360
X10050 1 2 DECAP7JI3V $T=205520 33600 1 180 $X=201170 $Y=32960
X10051 1 2 DECAP7JI3V $T=203280 42560 0 0 $X=202850 $Y=41920
X10052 1 2 DECAP7JI3V $T=215040 69440 1 0 $X=214610 $Y=64320
X10053 1 2 DECAP7JI3V $T=216160 60480 0 0 $X=215730 $Y=59840
X10054 1 2 DECAP7JI3V $T=218400 87360 1 0 $X=217970 $Y=82240
X10055 1 2 DECAP7JI3V $T=218960 69440 1 0 $X=218530 $Y=64320
X10056 1 2 DECAP7JI3V $T=220080 60480 0 0 $X=219650 $Y=59840
X10057 1 2 DECAP7JI3V $T=221200 33600 1 0 $X=220770 $Y=28480
X10058 1 2 DECAP7JI3V $T=221200 212800 0 0 $X=220770 $Y=212160
X10059 1 2 DECAP7JI3V $T=222320 24640 0 0 $X=221890 $Y=24000
X10060 1 2 DECAP7JI3V $T=222320 87360 1 0 $X=221890 $Y=82240
X10061 1 2 DECAP7JI3V $T=222880 69440 1 0 $X=222450 $Y=64320
X10062 1 2 DECAP7JI3V $T=222880 168000 0 0 $X=222450 $Y=167360
X10063 1 2 DECAP7JI3V $T=223440 185920 0 0 $X=223010 $Y=185280
X10064 1 2 DECAP7JI3V $T=224000 42560 0 0 $X=223570 $Y=41920
X10065 1 2 DECAP7JI3V $T=225120 33600 1 0 $X=224690 $Y=28480
X10066 1 2 DECAP7JI3V $T=225120 212800 0 0 $X=224690 $Y=212160
X10067 1 2 DECAP7JI3V $T=225680 212800 1 0 $X=225250 $Y=207680
X10068 1 2 DECAP7JI3V $T=226240 24640 0 0 $X=225810 $Y=24000
X10069 1 2 DECAP7JI3V $T=226240 87360 1 0 $X=225810 $Y=82240
X10070 1 2 DECAP7JI3V $T=226800 168000 0 0 $X=226370 $Y=167360
X10071 1 2 DECAP7JI3V $T=227360 185920 0 0 $X=226930 $Y=185280
X10072 1 2 DECAP7JI3V $T=227920 42560 0 0 $X=227490 $Y=41920
X10073 1 2 DECAP7JI3V $T=229040 78400 0 0 $X=228610 $Y=77760
X10074 1 2 DECAP7JI3V $T=229040 87360 0 0 $X=228610 $Y=86720
X10075 1 2 DECAP7JI3V $T=229040 96320 0 0 $X=228610 $Y=95680
X10076 1 2 DECAP7JI3V $T=229040 105280 0 0 $X=228610 $Y=104640
X10077 1 2 DECAP7JI3V $T=229040 132160 0 0 $X=228610 $Y=131520
X10078 1 2 DECAP7JI3V $T=231840 78400 1 0 $X=231410 $Y=73280
X10079 1 2 DECAP7JI3V $T=231840 123200 1 0 $X=231410 $Y=118080
X10080 1 2 DECAP7JI3V $T=232960 132160 0 0 $X=232530 $Y=131520
X10081 1 2 DECAP7JI3V $T=234080 141120 1 0 $X=233650 $Y=136000
X10082 1 2 DECAP7JI3V $T=235760 78400 1 0 $X=235330 $Y=73280
X10083 1 2 DECAP7JI3V $T=235760 123200 1 0 $X=235330 $Y=118080
X10084 1 2 DECAP7JI3V $T=239680 78400 1 0 $X=239250 $Y=73280
X10085 1 2 DECAP7JI3V $T=243600 78400 1 0 $X=243170 $Y=73280
X10086 1 2 DECAP7JI3V $T=249200 176960 0 180 $X=244850 $Y=171840
X10087 1 2 DECAP7JI3V $T=249200 176960 1 0 $X=248770 $Y=171840
X10088 1 2 DECAP7JI3V $T=251440 96320 1 0 $X=251010 $Y=91200
X10089 1 2 DECAP7JI3V $T=254240 185920 1 0 $X=253810 $Y=180800
X10090 1 2 DECAP7JI3V $T=258720 96320 0 0 $X=258290 $Y=95680
X10091 1 2 DECAP7JI3V $T=262640 96320 0 0 $X=262210 $Y=95680
X10092 1 2 DECAP7JI3V $T=266560 96320 0 0 $X=266130 $Y=95680
X10093 1 2 DECAP7JI3V $T=267120 78400 0 0 $X=266690 $Y=77760
X10094 1 2 DECAP7JI3V $T=267680 78400 1 0 $X=267250 $Y=73280
X10095 1 2 DECAP7JI3V $T=270480 24640 0 0 $X=270050 $Y=24000
X10096 1 2 DECAP7JI3V $T=270480 96320 0 0 $X=270050 $Y=95680
X10097 1 2 DECAP7JI3V $T=271040 78400 0 0 $X=270610 $Y=77760
X10098 1 2 DECAP7JI3V $T=271040 141120 1 0 $X=270610 $Y=136000
X10099 1 2 DECAP7JI3V $T=271040 141120 0 0 $X=270610 $Y=140480
X10100 1 2 DECAP7JI3V $T=271040 150080 1 0 $X=270610 $Y=144960
X10101 1 2 DECAP7JI3V $T=276640 203840 1 0 $X=276210 $Y=198720
X10102 1 2 DECAP7JI3V $T=280560 203840 1 0 $X=280130 $Y=198720
X10103 1 2 DECAP7JI3V $T=284480 203840 1 0 $X=284050 $Y=198720
X10104 1 2 DECAP7JI3V $T=285040 105280 1 0 $X=284610 $Y=100160
X10105 1 2 DECAP7JI3V $T=285600 185920 1 0 $X=285170 $Y=180800
X10106 1 2 DECAP7JI3V $T=288400 203840 1 0 $X=287970 $Y=198720
X10107 1 2 DECAP7JI3V $T=288960 105280 1 0 $X=288530 $Y=100160
X10108 1 2 DECAP7JI3V $T=291200 42560 1 0 $X=290770 $Y=37440
X10109 1 2 DECAP7JI3V $T=292320 132160 0 0 $X=291890 $Y=131520
X10110 1 2 DECAP7JI3V $T=297360 176960 0 0 $X=296930 $Y=176320
X10111 1 2 DECAP7JI3V $T=302960 96320 0 0 $X=302530 $Y=95680
X10112 1 2 DECAP7JI3V $T=306880 96320 0 0 $X=306450 $Y=95680
X10113 1 2 DECAP7JI3V $T=310240 159040 1 0 $X=309810 $Y=153920
X10114 1 2 DECAP7JI3V $T=310800 96320 0 0 $X=310370 $Y=95680
X10115 1 2 DECAP7JI3V $T=314720 78400 0 0 $X=314290 $Y=77760
X10116 1 2 DECAP7JI3V $T=316400 87360 0 0 $X=315970 $Y=86720
X10117 1 2 DECAP7JI3V $T=318640 141120 0 0 $X=318210 $Y=140480
X10118 1 2 DECAP7JI3V $T=320320 87360 0 0 $X=319890 $Y=86720
X10119 1 2 DECAP7JI3V $T=323120 194880 1 0 $X=322690 $Y=189760
X10120 1 2 DECAP7JI3V $T=324240 87360 0 0 $X=323810 $Y=86720
X10121 1 2 DECAP7JI3V $T=325360 123200 1 0 $X=324930 $Y=118080
X10122 1 2 DECAP7JI3V $T=326480 42560 0 0 $X=326050 $Y=41920
X10123 1 2 DECAP7JI3V $T=327040 194880 1 0 $X=326610 $Y=189760
X10124 1 2 DECAP7JI3V $T=329840 203840 1 0 $X=329410 $Y=198720
X10125 1 2 DECAP7JI3V $T=333760 60480 0 0 $X=333330 $Y=59840
X10126 1 2 DECAP7JI3V $T=337680 60480 0 0 $X=337250 $Y=59840
X10127 1 2 DECAP7JI3V $T=342720 51520 1 0 $X=342290 $Y=46400
X10128 1 2 DECAP7JI3V $T=343280 69440 1 0 $X=342850 $Y=64320
X10129 1 2 DECAP7JI3V $T=344400 78400 0 0 $X=343970 $Y=77760
X10130 1 2 DECAP7JI3V $T=344400 96320 0 0 $X=343970 $Y=95680
X10131 1 2 DECAP7JI3V $T=344960 168000 0 0 $X=344530 $Y=167360
X10132 1 2 DECAP7JI3V $T=345520 96320 1 0 $X=345090 $Y=91200
X10133 1 2 DECAP7JI3V $T=345520 114240 0 0 $X=345090 $Y=113600
X10134 1 2 DECAP7JI3V $T=347200 69440 1 0 $X=346770 $Y=64320
X10135 1 2 DECAP7JI3V $T=348320 51520 0 0 $X=347890 $Y=50880
X10136 1 2 DECAP7JI3V $T=348320 78400 0 0 $X=347890 $Y=77760
X10137 1 2 DECAP7JI3V $T=348320 96320 0 0 $X=347890 $Y=95680
X10138 1 2 DECAP7JI3V $T=349440 96320 1 0 $X=349010 $Y=91200
X10139 1 2 DECAP7JI3V $T=349440 114240 0 0 $X=349010 $Y=113600
X10140 1 2 DECAP7JI3V $T=349440 176960 1 0 $X=349010 $Y=171840
X10141 1 2 DECAP7JI3V $T=350000 33600 1 0 $X=349570 $Y=28480
X10142 1 2 DECAP7JI3V $T=351120 69440 1 0 $X=350690 $Y=64320
X10143 1 2 DECAP7JI3V $T=351680 168000 1 0 $X=351250 $Y=162880
X10144 1 2 DECAP7JI3V $T=351680 176960 0 0 $X=351250 $Y=176320
X10145 1 2 DECAP7JI3V $T=352240 60480 1 0 $X=351810 $Y=55360
X10146 1 2 DECAP7JI3V $T=352240 78400 0 0 $X=351810 $Y=77760
X10147 1 2 DECAP7JI3V $T=352240 87360 1 0 $X=351810 $Y=82240
X10148 1 2 DECAP7JI3V $T=352240 87360 0 0 $X=351810 $Y=86720
X10149 1 2 DECAP7JI3V $T=352240 96320 0 0 $X=351810 $Y=95680
X10150 1 2 DECAP7JI3V $T=352240 123200 1 0 $X=351810 $Y=118080
X10151 1 2 DECAP7JI3V $T=352240 123200 0 0 $X=351810 $Y=122560
X10152 1 2 DECAP7JI3V $T=352240 141120 0 0 $X=351810 $Y=140480
X10153 1 2 DECAP7JI3V $T=352240 159040 0 0 $X=351810 $Y=158400
X10154 1 2 DECAP7JI3V $T=353360 96320 1 0 $X=352930 $Y=91200
X10155 1 2 DECAP7JI3V $T=353360 114240 1 0 $X=352930 $Y=109120
X10156 1 2 DECAP7JI3V $T=353360 114240 0 0 $X=352930 $Y=113600
X10157 1 2 DECAP7JI3V $T=353360 176960 1 0 $X=352930 $Y=171840
X10158 1 2 DECAP7JI3V $T=353920 33600 1 0 $X=353490 $Y=28480
X10159 1 2 DECAP7JI3V $T=355040 132160 1 0 $X=354610 $Y=127040
X10160 1 2 DECAP7JI3V $T=355600 176960 0 0 $X=355170 $Y=176320
X10161 1 2 DECAP7JI3V $T=356160 60480 1 0 $X=355730 $Y=55360
X10162 1 2 DECAP7JI3V $T=356160 78400 0 0 $X=355730 $Y=77760
X10163 1 2 DECAP7JI3V $T=356160 87360 1 0 $X=355730 $Y=82240
X10164 1 2 DECAP7JI3V $T=356160 87360 0 0 $X=355730 $Y=86720
X10165 1 2 DECAP7JI3V $T=356160 96320 0 0 $X=355730 $Y=95680
X10166 1 2 DECAP7JI3V $T=356160 123200 1 0 $X=355730 $Y=118080
X10167 1 2 DECAP7JI3V $T=356160 123200 0 0 $X=355730 $Y=122560
X10168 1 2 DECAP7JI3V $T=357280 176960 1 0 $X=356850 $Y=171840
X10169 1 2 DECAP7JI3V $T=373520 168000 1 0 $X=373090 $Y=162880
X10170 1 2 DECAP7JI3V $T=376320 51520 0 0 $X=375890 $Y=50880
X10171 1 2 DECAP7JI3V $T=381360 114240 1 0 $X=380930 $Y=109120
X10172 1 2 DECAP7JI3V $T=382480 105280 1 0 $X=382050 $Y=100160
X10173 1 2 DECAP7JI3V $T=386400 105280 1 0 $X=385970 $Y=100160
X10174 1 2 DECAP7JI3V $T=388640 96320 1 0 $X=388210 $Y=91200
X10175 1 2 DECAP7JI3V $T=390320 105280 1 0 $X=389890 $Y=100160
X10176 1 2 DECAP7JI3V $T=394240 105280 1 0 $X=393810 $Y=100160
X10177 1 2 DECAP7JI3V $T=416640 33600 1 0 $X=416210 $Y=28480
X10178 1 2 DECAP7JI3V $T=416640 78400 1 0 $X=416210 $Y=73280
X10179 1 2 DECAP7JI3V $T=416640 96320 1 0 $X=416210 $Y=91200
X10180 1 2 DECAP7JI3V $T=416640 212800 0 0 $X=416210 $Y=212160
X10181 1 2 DECAP7JI3V $T=419440 114240 0 0 $X=419010 $Y=113600
X10182 1 2 DECAP7JI3V $T=419440 123200 0 0 $X=419010 $Y=122560
X10183 1 2 DECAP7JI3V $T=419440 159040 0 0 $X=419010 $Y=158400
X10184 1 2 DECAP7JI3V $T=420560 33600 1 0 $X=420130 $Y=28480
X10185 1 2 DECAP7JI3V $T=420560 78400 1 0 $X=420130 $Y=73280
X10186 1 2 DECAP7JI3V $T=420560 87360 1 0 $X=420130 $Y=82240
X10187 1 2 DECAP7JI3V $T=420560 96320 1 0 $X=420130 $Y=91200
X10188 1 2 DECAP7JI3V $T=420560 105280 0 0 $X=420130 $Y=104640
X10189 1 2 DECAP7JI3V $T=420560 114240 1 0 $X=420130 $Y=109120
X10190 1 2 DECAP7JI3V $T=420560 194880 1 0 $X=420130 $Y=189760
X10191 1 2 DECAP7JI3V $T=420560 212800 0 0 $X=420130 $Y=212160
X10192 1 2 DECAP7JI3V $T=423360 24640 0 0 $X=422930 $Y=24000
X10193 1 2 DECAP7JI3V $T=423360 114240 0 0 $X=422930 $Y=113600
X10194 1 2 DECAP7JI3V $T=423360 123200 0 0 $X=422930 $Y=122560
X10195 1 2 DECAP7JI3V $T=423360 159040 0 0 $X=422930 $Y=158400
X10196 1 2 DECAP7JI3V $T=423360 176960 1 0 $X=422930 $Y=171840
X10197 1 2 DECAP7JI3V $T=424480 33600 1 0 $X=424050 $Y=28480
X10198 1 2 DECAP7JI3V $T=424480 78400 1 0 $X=424050 $Y=73280
X10199 1 2 DECAP7JI3V $T=424480 87360 1 0 $X=424050 $Y=82240
X10200 1 2 DECAP7JI3V $T=424480 96320 1 0 $X=424050 $Y=91200
X10201 1 2 DECAP7JI3V $T=424480 105280 0 0 $X=424050 $Y=104640
X10202 1 2 DECAP7JI3V $T=424480 114240 1 0 $X=424050 $Y=109120
X10203 1 2 DECAP7JI3V $T=424480 123200 1 0 $X=424050 $Y=118080
X10204 1 2 DECAP7JI3V $T=424480 141120 1 0 $X=424050 $Y=136000
X10205 1 2 DECAP7JI3V $T=424480 194880 1 0 $X=424050 $Y=189760
X10206 1 2 DECAP7JI3V $T=424480 212800 0 0 $X=424050 $Y=212160
X10207 1 2 DECAP7JI3V $T=427280 24640 0 0 $X=426850 $Y=24000
X10208 1 2 DECAP7JI3V $T=427280 33600 0 0 $X=426850 $Y=32960
X10209 1 2 DECAP7JI3V $T=427280 42560 1 0 $X=426850 $Y=37440
X10210 1 2 DECAP7JI3V $T=427280 42560 0 0 $X=426850 $Y=41920
X10211 1 2 DECAP7JI3V $T=427280 51520 1 0 $X=426850 $Y=46400
X10212 1 2 DECAP7JI3V $T=427280 51520 0 0 $X=426850 $Y=50880
X10213 1 2 DECAP7JI3V $T=427280 60480 1 0 $X=426850 $Y=55360
X10214 1 2 DECAP7JI3V $T=427280 60480 0 0 $X=426850 $Y=59840
X10215 1 2 DECAP7JI3V $T=427280 69440 1 0 $X=426850 $Y=64320
X10216 1 2 DECAP7JI3V $T=427280 69440 0 0 $X=426850 $Y=68800
X10217 1 2 DECAP7JI3V $T=427280 87360 0 0 $X=426850 $Y=86720
X10218 1 2 DECAP7JI3V $T=427280 105280 1 0 $X=426850 $Y=100160
X10219 1 2 DECAP7JI3V $T=427280 114240 0 0 $X=426850 $Y=113600
X10220 1 2 DECAP7JI3V $T=427280 123200 0 0 $X=426850 $Y=122560
X10221 1 2 DECAP7JI3V $T=427280 159040 0 0 $X=426850 $Y=158400
X10222 1 2 DECAP7JI3V $T=427280 168000 0 0 $X=426850 $Y=167360
X10223 1 2 DECAP7JI3V $T=427280 176960 1 0 $X=426850 $Y=171840
X10224 1 2 DECAP7JI3V $T=427280 194880 0 0 $X=426850 $Y=194240
X10225 1 2 DECAP7JI3V $T=428400 24640 1 0 $X=427970 $Y=19520
X10226 1 2 DECAP7JI3V $T=428400 33600 1 0 $X=427970 $Y=28480
X10227 1 2 DECAP7JI3V $T=428400 78400 1 0 $X=427970 $Y=73280
X10228 1 2 DECAP7JI3V $T=428400 78400 0 0 $X=427970 $Y=77760
X10229 1 2 DECAP7JI3V $T=428400 87360 1 0 $X=427970 $Y=82240
X10230 1 2 DECAP7JI3V $T=428400 96320 1 0 $X=427970 $Y=91200
X10231 1 2 DECAP7JI3V $T=428400 96320 0 0 $X=427970 $Y=95680
X10232 1 2 DECAP7JI3V $T=428400 105280 0 0 $X=427970 $Y=104640
X10233 1 2 DECAP7JI3V $T=428400 114240 1 0 $X=427970 $Y=109120
X10234 1 2 DECAP7JI3V $T=428400 123200 1 0 $X=427970 $Y=118080
X10235 1 2 DECAP7JI3V $T=428400 141120 1 0 $X=427970 $Y=136000
X10236 1 2 DECAP7JI3V $T=428400 168000 1 0 $X=427970 $Y=162880
X10237 1 2 DECAP7JI3V $T=428400 194880 1 0 $X=427970 $Y=189760
X10238 1 2 DECAP7JI3V $T=428400 212800 1 0 $X=427970 $Y=207680
X10239 1 2 DECAP7JI3V $T=428400 212800 0 0 $X=427970 $Y=212160
X10240 1 2 DECAP7JI3V $T=431200 24640 0 0 $X=430770 $Y=24000
X10241 1 2 DECAP7JI3V $T=431200 33600 0 0 $X=430770 $Y=32960
X10242 1 2 DECAP7JI3V $T=431200 42560 1 0 $X=430770 $Y=37440
X10243 1 2 DECAP7JI3V $T=431200 42560 0 0 $X=430770 $Y=41920
X10244 1 2 DECAP7JI3V $T=431200 51520 1 0 $X=430770 $Y=46400
X10245 1 2 DECAP7JI3V $T=431200 51520 0 0 $X=430770 $Y=50880
X10246 1 2 DECAP7JI3V $T=431200 60480 1 0 $X=430770 $Y=55360
X10247 1 2 DECAP7JI3V $T=431200 60480 0 0 $X=430770 $Y=59840
X10248 1 2 DECAP7JI3V $T=431200 69440 1 0 $X=430770 $Y=64320
X10249 1 2 DECAP7JI3V $T=431200 69440 0 0 $X=430770 $Y=68800
X10250 1 2 DECAP7JI3V $T=431200 87360 0 0 $X=430770 $Y=86720
X10251 1 2 DECAP7JI3V $T=431200 105280 1 0 $X=430770 $Y=100160
X10252 1 2 DECAP7JI3V $T=431200 114240 0 0 $X=430770 $Y=113600
X10253 1 2 DECAP7JI3V $T=431200 123200 0 0 $X=430770 $Y=122560
X10254 1 2 DECAP7JI3V $T=431200 150080 0 0 $X=430770 $Y=149440
X10255 1 2 DECAP7JI3V $T=431200 159040 0 0 $X=430770 $Y=158400
X10256 1 2 DECAP7JI3V $T=431200 168000 0 0 $X=430770 $Y=167360
X10257 1 2 DECAP7JI3V $T=431200 176960 1 0 $X=430770 $Y=171840
X10258 1 2 DECAP7JI3V $T=431200 176960 0 0 $X=430770 $Y=176320
X10259 1 2 DECAP7JI3V $T=431200 185920 1 0 $X=430770 $Y=180800
X10260 1 2 DECAP7JI3V $T=431200 194880 0 0 $X=430770 $Y=194240
X10261 1 2 DECAP7JI3V $T=431200 203840 1 0 $X=430770 $Y=198720
X10262 1 2 DECAP5JI3V $T=20160 105280 0 0 $X=19730 $Y=104640
X10263 1 2 DECAP5JI3V $T=20160 114240 1 0 $X=19730 $Y=109120
X10264 1 2 DECAP5JI3V $T=20160 123200 0 0 $X=19730 $Y=122560
X10265 1 2 DECAP5JI3V $T=20160 132160 1 0 $X=19730 $Y=127040
X10266 1 2 DECAP5JI3V $T=20160 132160 0 0 $X=19730 $Y=131520
X10267 1 2 DECAP5JI3V $T=20160 194880 1 0 $X=19730 $Y=189760
X10268 1 2 DECAP5JI3V $T=36960 114240 0 0 $X=36530 $Y=113600
X10269 1 2 DECAP5JI3V $T=42000 42560 1 0 $X=41570 $Y=37440
X10270 1 2 DECAP5JI3V $T=42000 42560 0 0 $X=41570 $Y=41920
X10271 1 2 DECAP5JI3V $T=42000 51520 1 0 $X=41570 $Y=46400
X10272 1 2 DECAP5JI3V $T=42000 51520 0 0 $X=41570 $Y=50880
X10273 1 2 DECAP5JI3V $T=42560 60480 1 0 $X=42130 $Y=55360
X10274 1 2 DECAP5JI3V $T=48160 176960 1 0 $X=47730 $Y=171840
X10275 1 2 DECAP5JI3V $T=48160 203840 1 0 $X=47730 $Y=198720
X10276 1 2 DECAP5JI3V $T=54320 24640 1 0 $X=53890 $Y=19520
X10277 1 2 DECAP5JI3V $T=59920 42560 1 0 $X=59490 $Y=37440
X10278 1 2 DECAP5JI3V $T=60480 60480 0 0 $X=60050 $Y=59840
X10279 1 2 DECAP5JI3V $T=62160 78400 0 0 $X=61730 $Y=77760
X10280 1 2 DECAP5JI3V $T=62160 87360 0 0 $X=61730 $Y=86720
X10281 1 2 DECAP5JI3V $T=62720 105280 0 0 $X=62290 $Y=104640
X10282 1 2 DECAP5JI3V $T=63280 114240 0 0 $X=62850 $Y=113600
X10283 1 2 DECAP5JI3V $T=67760 159040 1 0 $X=67330 $Y=153920
X10284 1 2 DECAP5JI3V $T=72240 212800 1 0 $X=71810 $Y=207680
X10285 1 2 DECAP5JI3V $T=94080 51520 1 0 $X=93650 $Y=46400
X10286 1 2 DECAP5JI3V $T=94080 51520 0 0 $X=93650 $Y=50880
X10287 1 2 DECAP5JI3V $T=94080 60480 1 0 $X=93650 $Y=55360
X10288 1 2 DECAP5JI3V $T=95760 150080 1 0 $X=95330 $Y=144960
X10289 1 2 DECAP5JI3V $T=98560 185920 1 0 $X=98130 $Y=180800
X10290 1 2 DECAP5JI3V $T=100240 105280 1 0 $X=99810 $Y=100160
X10291 1 2 DECAP5JI3V $T=100240 123200 0 0 $X=99810 $Y=122560
X10292 1 2 DECAP5JI3V $T=100240 132160 1 0 $X=99810 $Y=127040
X10293 1 2 DECAP5JI3V $T=100240 141120 0 0 $X=99810 $Y=140480
X10294 1 2 DECAP5JI3V $T=100240 159040 1 0 $X=99810 $Y=153920
X10295 1 2 DECAP5JI3V $T=107520 105280 0 0 $X=107090 $Y=104640
X10296 1 2 DECAP5JI3V $T=108080 87360 0 0 $X=107650 $Y=86720
X10297 1 2 DECAP5JI3V $T=108640 78400 0 0 $X=108210 $Y=77760
X10298 1 2 DECAP5JI3V $T=110880 114240 1 0 $X=110450 $Y=109120
X10299 1 2 DECAP5JI3V $T=115360 114240 0 0 $X=114930 $Y=113600
X10300 1 2 DECAP5JI3V $T=121520 24640 1 180 $X=118290 $Y=24000
X10301 1 2 DECAP5JI3V $T=119280 168000 0 0 $X=118850 $Y=167360
X10302 1 2 DECAP5JI3V $T=134960 24640 1 0 $X=134530 $Y=19520
X10303 1 2 DECAP5JI3V $T=140000 78400 0 0 $X=139570 $Y=77760
X10304 1 2 DECAP5JI3V $T=140000 87360 0 0 $X=139570 $Y=86720
X10305 1 2 DECAP5JI3V $T=142800 69440 0 0 $X=142370 $Y=68800
X10306 1 2 DECAP5JI3V $T=156240 212800 0 0 $X=155810 $Y=212160
X10307 1 2 DECAP5JI3V $T=159600 78400 1 0 $X=159170 $Y=73280
X10308 1 2 DECAP5JI3V $T=163520 168000 1 0 $X=163090 $Y=162880
X10309 1 2 DECAP5JI3V $T=166320 33600 0 0 $X=165890 $Y=32960
X10310 1 2 DECAP5JI3V $T=179760 60480 1 0 $X=179330 $Y=55360
X10311 1 2 DECAP5JI3V $T=181440 168000 1 0 $X=181010 $Y=162880
X10312 1 2 DECAP5JI3V $T=184240 87360 1 0 $X=183810 $Y=82240
X10313 1 2 DECAP5JI3V $T=184800 42560 1 0 $X=184370 $Y=37440
X10314 1 2 DECAP5JI3V $T=185360 132160 1 0 $X=184930 $Y=127040
X10315 1 2 DECAP5JI3V $T=188720 212800 1 0 $X=188290 $Y=207680
X10316 1 2 DECAP5JI3V $T=197680 51520 1 0 $X=197250 $Y=46400
X10317 1 2 DECAP5JI3V $T=197680 51520 0 0 $X=197250 $Y=50880
X10318 1 2 DECAP5JI3V $T=224000 51520 1 0 $X=223570 $Y=46400
X10319 1 2 DECAP5JI3V $T=224000 60480 0 0 $X=223570 $Y=59840
X10320 1 2 DECAP5JI3V $T=224000 176960 0 0 $X=223570 $Y=176320
X10321 1 2 DECAP5JI3V $T=224000 185920 1 0 $X=223570 $Y=180800
X10322 1 2 DECAP5JI3V $T=228480 141120 0 0 $X=228050 $Y=140480
X10323 1 2 DECAP5JI3V $T=228480 150080 0 0 $X=228050 $Y=149440
X10324 1 2 DECAP5JI3V $T=229040 33600 1 0 $X=228610 $Y=28480
X10325 1 2 DECAP5JI3V $T=229040 212800 0 0 $X=228610 $Y=212160
X10326 1 2 DECAP5JI3V $T=230160 24640 0 0 $X=229730 $Y=24000
X10327 1 2 DECAP5JI3V $T=230160 87360 1 0 $X=229730 $Y=82240
X10328 1 2 DECAP5JI3V $T=230720 168000 0 0 $X=230290 $Y=167360
X10329 1 2 DECAP5JI3V $T=231840 114240 1 0 $X=231410 $Y=109120
X10330 1 2 DECAP5JI3V $T=237440 123200 0 0 $X=237010 $Y=122560
X10331 1 2 DECAP5JI3V $T=244160 33600 1 0 $X=243730 $Y=28480
X10332 1 2 DECAP5JI3V $T=251440 114240 1 0 $X=251010 $Y=109120
X10333 1 2 DECAP5JI3V $T=263760 176960 1 0 $X=263330 $Y=171840
X10334 1 2 DECAP5JI3V $T=272160 132160 1 0 $X=271730 $Y=127040
X10335 1 2 DECAP5JI3V $T=273280 60480 1 0 $X=272850 $Y=55360
X10336 1 2 DECAP5JI3V $T=274400 123200 0 0 $X=273970 $Y=122560
X10337 1 2 DECAP5JI3V $T=276080 203840 0 0 $X=275650 $Y=203200
X10338 1 2 DECAP5JI3V $T=277760 132160 0 0 $X=277330 $Y=131520
X10339 1 2 DECAP5JI3V $T=278320 33600 0 0 $X=277890 $Y=32960
X10340 1 2 DECAP5JI3V $T=285040 33600 1 0 $X=284610 $Y=28480
X10341 1 2 DECAP5JI3V $T=285600 114240 0 0 $X=285170 $Y=113600
X10342 1 2 DECAP5JI3V $T=294000 51520 0 180 $X=290770 $Y=46400
X10343 1 2 DECAP5JI3V $T=291200 51520 0 0 $X=290770 $Y=50880
X10344 1 2 DECAP5JI3V $T=291200 60480 1 0 $X=290770 $Y=55360
X10345 1 2 DECAP5JI3V $T=291200 60480 0 0 $X=290770 $Y=59840
X10346 1 2 DECAP5JI3V $T=291760 96320 1 0 $X=291330 $Y=91200
X10347 1 2 DECAP5JI3V $T=299040 159040 1 0 $X=298610 $Y=153920
X10348 1 2 DECAP5JI3V $T=301840 33600 0 0 $X=301410 $Y=32960
X10349 1 2 DECAP5JI3V $T=306880 194880 1 0 $X=306450 $Y=189760
X10350 1 2 DECAP5JI3V $T=309120 60480 0 0 $X=308690 $Y=59840
X10351 1 2 DECAP5JI3V $T=312480 212800 1 0 $X=312050 $Y=207680
X10352 1 2 DECAP5JI3V $T=314160 114240 0 0 $X=313730 $Y=113600
X10353 1 2 DECAP5JI3V $T=317520 24640 0 0 $X=317090 $Y=24000
X10354 1 2 DECAP5JI3V $T=327040 78400 1 0 $X=326610 $Y=73280
X10355 1 2 DECAP5JI3V $T=327040 194880 0 0 $X=326610 $Y=194240
X10356 1 2 DECAP5JI3V $T=328720 69440 0 0 $X=328290 $Y=68800
X10357 1 2 DECAP5JI3V $T=342720 212800 1 0 $X=342290 $Y=207680
X10358 1 2 DECAP5JI3V $T=352240 51520 0 0 $X=351810 $Y=50880
X10359 1 2 DECAP5JI3V $T=355040 159040 1 0 $X=354610 $Y=153920
X10360 1 2 DECAP5JI3V $T=355600 141120 1 0 $X=355170 $Y=136000
X10361 1 2 DECAP5JI3V $T=355600 150080 1 0 $X=355170 $Y=144960
X10362 1 2 DECAP5JI3V $T=355600 168000 1 0 $X=355170 $Y=162880
X10363 1 2 DECAP5JI3V $T=357280 96320 1 0 $X=356850 $Y=91200
X10364 1 2 DECAP5JI3V $T=357280 114240 0 0 $X=356850 $Y=113600
X10365 1 2 DECAP5JI3V $T=357840 33600 1 0 $X=357410 $Y=28480
X10366 1 2 DECAP5JI3V $T=358400 105280 1 0 $X=357970 $Y=100160
X10367 1 2 DECAP5JI3V $T=362880 51520 0 180 $X=359650 $Y=46400
X10368 1 2 DECAP5JI3V $T=360080 60480 1 0 $X=359650 $Y=55360
X10369 1 2 DECAP5JI3V $T=377440 60480 0 0 $X=377010 $Y=59840
X10370 1 2 DECAP5JI3V $T=383040 132160 0 180 $X=379810 $Y=127040
X10371 1 2 DECAP5JI3V $T=381360 105280 0 0 $X=380930 $Y=104640
X10372 1 2 DECAP5JI3V $T=381360 123200 1 0 $X=380930 $Y=118080
X10373 1 2 DECAP5JI3V $T=381920 114240 0 0 $X=381490 $Y=113600
X10374 1 2 DECAP5JI3V $T=381920 141120 0 0 $X=381490 $Y=140480
X10375 1 2 DECAP5JI3V $T=385840 33600 1 0 $X=385410 $Y=28480
X10376 1 2 DECAP5JI3V $T=393680 150080 1 180 $X=390450 $Y=149440
X10377 1 2 DECAP5JI3V $T=392560 96320 1 0 $X=392130 $Y=91200
X10378 1 2 DECAP5JI3V $T=395360 42560 1 0 $X=394930 $Y=37440
X10379 1 2 DECAP5JI3V $T=395360 42560 0 0 $X=394930 $Y=41920
X10380 1 2 DECAP5JI3V $T=395360 60480 1 0 $X=394930 $Y=55360
X10381 1 2 DECAP5JI3V $T=395360 60480 0 0 $X=394930 $Y=59840
X10382 1 2 DECAP5JI3V $T=395360 69440 1 0 $X=394930 $Y=64320
X10383 1 2 DECAP5JI3V $T=395360 69440 0 0 $X=394930 $Y=68800
X10384 1 2 DECAP5JI3V $T=409360 24640 1 180 $X=406130 $Y=24000
X10385 1 2 DECAP5JI3V $T=432320 24640 1 0 $X=431890 $Y=19520
X10386 1 2 DECAP5JI3V $T=432320 33600 1 0 $X=431890 $Y=28480
X10387 1 2 DECAP5JI3V $T=432320 78400 1 0 $X=431890 $Y=73280
X10388 1 2 DECAP5JI3V $T=432320 78400 0 0 $X=431890 $Y=77760
X10389 1 2 DECAP5JI3V $T=432320 87360 1 0 $X=431890 $Y=82240
X10390 1 2 DECAP5JI3V $T=432320 96320 1 0 $X=431890 $Y=91200
X10391 1 2 DECAP5JI3V $T=432320 96320 0 0 $X=431890 $Y=95680
X10392 1 2 DECAP5JI3V $T=432320 105280 0 0 $X=431890 $Y=104640
X10393 1 2 DECAP5JI3V $T=432320 114240 1 0 $X=431890 $Y=109120
X10394 1 2 DECAP5JI3V $T=432320 123200 1 0 $X=431890 $Y=118080
X10395 1 2 DECAP5JI3V $T=432320 132160 1 0 $X=431890 $Y=127040
X10396 1 2 DECAP5JI3V $T=432320 141120 1 0 $X=431890 $Y=136000
X10397 1 2 DECAP5JI3V $T=432320 159040 1 0 $X=431890 $Y=153920
X10398 1 2 DECAP5JI3V $T=432320 168000 1 0 $X=431890 $Y=162880
X10399 1 2 DECAP5JI3V $T=432320 194880 1 0 $X=431890 $Y=189760
X10400 1 2 DECAP5JI3V $T=432320 212800 1 0 $X=431890 $Y=207680
X10401 1 2 DECAP5JI3V $T=432320 212800 0 0 $X=431890 $Y=212160
X10402 1 2 DECAP10JI3V $T=20160 114240 0 0 $X=19730 $Y=113600
X10403 1 2 DECAP10JI3V $T=20160 123200 1 0 $X=19730 $Y=118080
X10404 1 2 DECAP10JI3V $T=20160 159040 1 0 $X=19730 $Y=153920
X10405 1 2 DECAP10JI3V $T=20160 176960 0 0 $X=19730 $Y=176320
X10406 1 2 DECAP10JI3V $T=20160 185920 0 0 $X=19730 $Y=185280
X10407 1 2 DECAP10JI3V $T=34160 24640 0 0 $X=33730 $Y=24000
X10408 1 2 DECAP10JI3V $T=34160 87360 1 0 $X=33730 $Y=82240
X10409 1 2 DECAP10JI3V $T=34160 194880 0 0 $X=33730 $Y=194240
X10410 1 2 DECAP10JI3V $T=39760 123200 0 0 $X=39330 $Y=122560
X10411 1 2 DECAP10JI3V $T=76160 203840 1 0 $X=75730 $Y=198720
X10412 1 2 DECAP10JI3V $T=77840 141120 0 0 $X=77410 $Y=140480
X10413 1 2 DECAP10JI3V $T=90720 176960 1 0 $X=90290 $Y=171840
X10414 1 2 DECAP10JI3V $T=92960 168000 0 0 $X=92530 $Y=167360
X10415 1 2 DECAP10JI3V $T=95200 159040 0 0 $X=94770 $Y=158400
X10416 1 2 DECAP10JI3V $T=95760 176960 0 0 $X=95330 $Y=176320
X10417 1 2 DECAP10JI3V $T=100240 194880 1 0 $X=99810 $Y=189760
X10418 1 2 DECAP10JI3V $T=140560 176960 1 0 $X=140130 $Y=171840
X10419 1 2 DECAP10JI3V $T=151760 132160 0 0 $X=151330 $Y=131520
X10420 1 2 DECAP10JI3V $T=152880 87360 1 0 $X=152450 $Y=82240
X10421 1 2 DECAP10JI3V $T=204400 123200 1 0 $X=203970 $Y=118080
X10422 1 2 DECAP10JI3V $T=212240 42560 1 0 $X=211810 $Y=37440
X10423 1 2 DECAP10JI3V $T=221200 51520 0 0 $X=220770 $Y=50880
X10424 1 2 DECAP10JI3V $T=223440 78400 0 0 $X=223010 $Y=77760
X10425 1 2 DECAP10JI3V $T=223440 87360 0 0 $X=223010 $Y=86720
X10426 1 2 DECAP10JI3V $T=223440 96320 0 0 $X=223010 $Y=95680
X10427 1 2 DECAP10JI3V $T=223440 105280 0 0 $X=223010 $Y=104640
X10428 1 2 DECAP10JI3V $T=223440 132160 0 0 $X=223010 $Y=131520
X10429 1 2 DECAP10JI3V $T=223440 159040 1 0 $X=223010 $Y=153920
X10430 1 2 DECAP10JI3V $T=224560 176960 1 0 $X=224130 $Y=171840
X10431 1 2 DECAP10JI3V $T=226240 123200 1 0 $X=225810 $Y=118080
X10432 1 2 DECAP10JI3V $T=228480 141120 1 0 $X=228050 $Y=136000
X10433 1 2 DECAP10JI3V $T=243040 150080 1 0 $X=242610 $Y=144960
X10434 1 2 DECAP10JI3V $T=245840 96320 1 0 $X=245410 $Y=91200
X10435 1 2 DECAP10JI3V $T=253120 105280 0 0 $X=252690 $Y=104640
X10436 1 2 DECAP10JI3V $T=283360 150080 0 0 $X=282930 $Y=149440
X10437 1 2 DECAP10JI3V $T=285600 42560 1 0 $X=285170 $Y=37440
X10438 1 2 DECAP10JI3V $T=308560 176960 0 0 $X=308130 $Y=176320
X10439 1 2 DECAP10JI3V $T=309120 78400 0 0 $X=308690 $Y=77760
X10440 1 2 DECAP10JI3V $T=318640 123200 1 0 $X=318210 $Y=118080
X10441 1 2 DECAP10JI3V $T=326480 105280 0 0 $X=326050 $Y=104640
X10442 1 2 DECAP10JI3V $T=338800 78400 0 0 $X=338370 $Y=77760
X10443 1 2 DECAP10JI3V $T=340480 33600 1 0 $X=340050 $Y=28480
X10444 1 2 DECAP10JI3V $T=347760 114240 1 0 $X=347330 $Y=109120
X10445 1 2 DECAP10JI3V $T=352240 42560 1 0 $X=351810 $Y=37440
X10446 1 2 DECAP10JI3V $T=352240 105280 0 0 $X=351810 $Y=104640
X10447 1 2 DECAP10JI3V $T=352240 185920 0 0 $X=351810 $Y=185280
X10448 1 2 DECAP10JI3V $T=352800 168000 0 0 $X=352370 $Y=167360
X10449 1 2 DECAP10JI3V $T=356720 42560 0 0 $X=356290 $Y=41920
X10450 1 2 DECAP10JI3V $T=356720 60480 0 0 $X=356290 $Y=59840
X10451 1 2 DECAP10JI3V $T=373520 185920 0 180 $X=367490 $Y=180800
X10452 1 2 DECAP10JI3V $T=371280 69440 1 0 $X=370850 $Y=64320
X10453 1 2 DECAP10JI3V $T=413840 123200 0 0 $X=413410 $Y=122560
X10454 1 2 DECAP10JI3V $T=413840 159040 0 0 $X=413410 $Y=158400
X10455 1 2 DECAP10JI3V $T=421680 33600 0 0 $X=421250 $Y=32960
X10456 1 2 DECAP10JI3V $T=421680 60480 1 0 $X=421250 $Y=55360
X10457 1 2 DECAP10JI3V $T=421680 87360 0 0 $X=421250 $Y=86720
X10458 1 2 DECAP10JI3V $T=421680 168000 0 0 $X=421250 $Y=167360
D0 83 1 p_ddnwmv AREA=8.49716e-08 PJ=0.00124444 perimeter=0.00124444 $X=17730 $Y=17520 $dt=2
D1 2 1 p_dipdnwmv AREA=1.68269e-09 PJ=0.000846738 perimeter=0.000846738 $X=24380 $Y=192640 $dt=3
D2 2 1 p_dipdnwmv AREA=1.71436e-09 PJ=0.000856626 perimeter=0.000856626 $X=29010 $Y=138870 $dt=3
D3 2 1 p_dipdnwmv AREA=1.70244e-09 PJ=0.00085168 perimeter=0.00085168 $X=30130 $Y=120950 $dt=3
D4 2 1 p_dipdnwmv AREA=1.7101e-09 PJ=0.000852491 perimeter=0.000852491 $X=46940 $Y=94080 $dt=3
D5 2 1 p_dipdnwmv AREA=1.72326e-09 PJ=0.000856437 perimeter=0.000856437 $X=69890 $Y=67190 $dt=3
D6 2 1 p_dipdnwmv AREA=1.68194e-09 PJ=0.000847719 perimeter=0.000847719 $X=76460 $Y=210560 $dt=3
D7 2 1 p_dipdnwmv AREA=1.72011e-09 PJ=0.000854508 perimeter=0.000854508 $X=85570 $Y=85110 $dt=3
D8 2 1 p_dipdnwmv AREA=1.68085e-09 PJ=0.000847368 perimeter=0.000847368 $X=85570 $Y=201590 $dt=3
D9 2 1 p_dipdnwmv AREA=1.67889e-09 PJ=0.000849321 perimeter=0.000849321 $X=87810 $Y=165750 $dt=3
D10 2 1 p_dipdnwmv AREA=1.7123e-09 PJ=0.000855368 perimeter=0.000855368 $X=89490 $Y=147830 $dt=3
D11 2 1 p_dipdnwmv AREA=1.66499e-09 PJ=0.000851237 perimeter=0.000851237 $X=117490 $Y=31350 $dt=3
D12 2 1 p_dipdnwmv AREA=1.71216e-09 PJ=0.000861885 perimeter=0.000861885 $X=129810 $Y=40310 $dt=3
D13 2 1 p_dipdnwmv AREA=1.67656e-09 PJ=0.000846569 perimeter=0.000846569 $X=132610 $Y=183670 $dt=3
D14 2 1 p_dipdnwmv AREA=1.72262e-09 PJ=0.000856557 perimeter=0.000856557 $X=146610 $Y=58230 $dt=3
D15 2 1 p_dipdnwmv AREA=1.70024e-09 PJ=0.000851249 perimeter=0.000851249 $X=167890 $Y=111990 $dt=3
D16 2 1 p_dipdnwmv AREA=1.71539e-09 PJ=0.000856066 perimeter=0.000856066 $X=175170 $Y=129910 $dt=3
D17 2 1 p_dipdnwmv AREA=1.71256e-09 PJ=0.000853309 perimeter=0.000853309 $X=191410 $Y=103030 $dt=3
D18 2 1 p_dipdnwmv AREA=1.69697e-09 PJ=0.000852039 perimeter=0.000852039 $X=293890 $Y=156790 $dt=3
D19 2 1 p_dipdnwmv AREA=1.67952e-09 PJ=0.000847075 perimeter=0.000847075 $X=344380 $Y=174710 $dt=3
D20 2 1 p_dipdnwmv AREA=1.64744e-09 PJ=0.0008401 perimeter=0.0008401 $X=386290 $Y=22390 $dt=3
D21 2 1 p_dipdnwmv AREA=1.71423e-09 PJ=0.000853703 perimeter=0.000853703 $X=390210 $Y=76150 $dt=3
D22 2 1 p_dipdnwmv AREA=1.72604e-09 PJ=0.000856428 perimeter=0.000856428 $X=413730 $Y=49270 $dt=3
.ends aska_dig

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: aska_dig_lvs                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt aska_dig_lvs gndd vdd3
** N=83 EP=2 FDC=26952
X0 vdd3 gndd 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70
+ 71 72 73 74 75 76 77 78 79 80
+ 81 82 aska_dig $T=14565 6815 0 0 $X=14645 $Y=6815
.ends aska_dig_lvs
