* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : aska_dig_lvs                                 *
* Netlisted  : Mon Jul 15 19:51:23 2024                     *
* PVS Version: 23.10-p043 Mon Oct 2 18:09:08 PDT 2023      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(ne3i) nemi ndiff(D) p1trm(G) ndiff(S) pwitrm(B)
*.DEVTMPLT 1 MP(pe3i) pemi pdiff(D) p1trm(G) pdiff(S) dnwtrm(B)
*.DEVTMPLT 2 D(p_ddnwmv) p_ddnwmv bulk(POS) dnwtrm(NEG)
*.DEVTMPLT 3 D(p_dipdnwmv) p_dipwmv pwitrm(POS) dnwtrm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX2                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX2 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=6
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=6e-07 AD=2.96727e-13 AS=2.88e-13 PD=1.69091e-06 PS=2.16e-06 $X=620 $Y=950 $dt=0
M1 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=7.2e-07 AD=2.016e-13 AS=3.56073e-13 PD=1.512e-06 PS=2.02909e-06 $X=1590 $Y=830 $dt=0
M2 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=4.648e-13 AS=1.344e-13 PD=3.52e-06 PS=1.008e-06 $X=2480 $Y=1070 $dt=0
M3 vdd3i! A 6 vdd3i! pe3i L=3e-07 W=1.1e-06 AD=5.39943e-13 AS=5.28e-13 PD=2.20442e-06 PS=3.16e-06 $X=620 $Y=2410 $dt=1
M4 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=7.16507e-13 PD=1.87971e-06 PS=2.92528e-06 $X=1640 $Y=2410 $dt=1
M5 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=8.6265e-13 AS=2.751e-13 PD=4.56971e-06 PS=1.87971e-06 $X=2480 $Y=2410 $dt=1
.ends BUJI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND2JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND2JI3VX1 vdd3i! gnd3i! A B Q
*.DEVICECLIMB
** N=8 EP=5 FDC=6
M0 7 A 8 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=2.688e-13 PD=8.1e-07 PS=2.08e-06 $X=820 $Y=990 $dt=0
M1 gnd3i! B 7 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=2.57137e-13 AS=7e-14 PD=1.43669e-06 PS=8.1e-07 $X=1420 $Y=990 $dt=0
M2 Q 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=4.08663e-13 PD=2.74e-06 PS=2.28331e-06 $X=2390 $Y=660 $dt=0
M3 8 A vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=7.276e-13 PD=1.24e-06 PS=4.56e-06 $X=580 $Y=2410 $dt=1
M4 vdd3i! B 8 vdd3i! pe3i L=3e-07 W=7e-07 AD=3.64829e-13 AS=1.89e-13 PD=1.6455e-06 PS=1.24e-06 $X=1420 $Y=2410 $dt=1
M5 Q 8 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=7.34871e-13 PD=3.78e-06 PS=3.3145e-06 $X=2440 $Y=2410 $dt=1
.ends AND2JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: EN2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt EN2JI3VX0 vdd3i! gnd3i! A B Q
*.DEVICECLIMB
** N=10 EP=5 FDC=10
M0 8 A 9 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=620 $Y=980 $dt=0
M1 gnd3i! B 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=1220 $Y=980 $dt=0
M2 7 A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=1.134e-13 PD=9.6e-07 PS=9.6e-07 $X=2110 $Y=980 $dt=0
M3 gnd3i! B 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.698e-13 AS=1.134e-13 PD=3.22e-06 PS=9.6e-07 $X=3000 $Y=980 $dt=0
M4 Q 9 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=2.058e-13 PD=1.8e-06 PS=1.82e-06 $X=4440 $Y=1020 $dt=0
M5 9 A vdd3i! vdd3i! pe3i L=3e-07 W=9e-07 AD=3.195e-13 AS=8.517e-13 PD=1.61e-06 PS=4.61e-06 $X=685 $Y=2410 $dt=1
M6 vdd3i! B 9 vdd3i! pe3i L=3e-07 W=9e-07 AD=4.30855e-13 AS=3.195e-13 PD=1.83273e-06 PS=1.61e-06 $X=1695 $Y=2410 $dt=1
M7 10 A vdd3i! vdd3i! pe3i L=3e-07 W=1.3e-06 AD=1.95e-13 AS=6.22345e-13 PD=1.6e-06 PS=2.64727e-06 $X=2825 $Y=2520 $dt=1
M8 Q B 10 vdd3i! pe3i L=3e-07 W=1.3e-06 AD=6.21324e-13 AS=1.95e-13 PD=2.52941e-06 PS=1.6e-06 $X=3425 $Y=2520 $dt=1
M9 vdd3i! 9 Q vdd3i! pe3i L=3e-07 W=9.1e-07 AD=8.0675e-13 AS=4.34926e-13 PD=4.39e-06 PS=1.77059e-06 $X=4575 $Y=2520 $dt=1
.ends EN2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA2I1JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA2I1JI3VX1 vdd3i! gnd3i! AN Q B
*.DEVICECLIMB
** N=8 EP=5 FDC=6
M0 gnd3i! AN 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.44754e-13 AS=2.016e-13 PD=1.25038e-06 PS=1.8e-06 $X=620 $Y=660 $dt=0
M1 7 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=5.18646e-13 PD=1.14e-06 PS=2.64962e-06 $X=1680 $Y=660 $dt=0
M2 Q B 7 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=1.1125e-13 PD=2.74e-06 PS=1.14e-06 $X=2280 $Y=660 $dt=0
M3 vdd3i! AN 8 vdd3i! pe3i L=3e-07 W=7e-07 AD=6.84341e-13 AS=3.36e-13 PD=3.08e-06 PS=2.36e-06 $X=620 $Y=2410 $dt=1
M4 Q 8 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.7e-13 AS=9.7763e-13 PD=1.54e-06 PS=4.4e-06 $X=1510 $Y=2410 $dt=1
M5 vdd3i! B Q vdd3i! pe3i L=3e-07 W=1e-06 AD=9.7763e-13 AS=2.7e-13 PD=4.4e-06 PS=1.54e-06 $X=2350 $Y=2410 $dt=1
.ends NA2I1JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO3I2JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO3I2JI3VX1 vdd3i! gnd3i! AN BN C Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 8 AN 9 gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=6e-14 AS=2.304e-13 PD=7.3e-07 PS=1.92e-06 $X=620 $Y=1070 $dt=0
M1 gnd3i! BN 8 gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=1.98937e-13 AS=6e-14 PD=1.31617e-06 PS=7.3e-07 $X=1220 $Y=1070 $dt=0
M2 Q C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.68863e-13 PD=1.43e-06 PS=2.4404e-06 $X=2060 $Y=660 $dt=0
M3 gnd3i! 9 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.329e-13 AS=2.403e-13 PD=2.77e-06 PS=1.43e-06 $X=2950 $Y=660 $dt=0
M4 9 AN vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=5.71409e-13 PD=1.24e-06 PS=2.5758e-06 $X=560 $Y=2590 $dt=1
M5 vdd3i! BN 9 vdd3i! pe3i L=3e-07 W=7e-07 AD=5.71409e-13 AS=1.89e-13 PD=2.5758e-06 PS=1.24e-06 $X=1400 $Y=2590 $dt=1
M6 10 C vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=1.15098e-12 PD=1.66e-06 PS=5.1884e-06 $X=2330 $Y=2410 $dt=1
M7 Q 9 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=8.46e-13 AS=1.7625e-13 PD=4.02e-06 PS=1.66e-06 $X=2880 $Y=2410 $dt=1
.ends NO3I2JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA2JI3VX1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA2JI3VX1 vdd3i! gnd3i! B Q A
*.DEVICECLIMB
** N=7 EP=5 FDC=4
M0 7 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=6.222e-13 PD=1.14e-06 PS=3.54e-06 $X=670 $Y=660 $dt=0
M1 Q A 7 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=1.1125e-13 PD=2.74e-06 PS=1.14e-06 $X=1270 $Y=660 $dt=0
M2 Q B vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.7e-13 AS=9.404e-13 PD=1.54e-06 PS=5.24e-06 $X=550 $Y=2410 $dt=1
M3 vdd3i! A Q vdd3i! pe3i L=3e-07 W=1e-06 AD=9.404e-13 AS=2.7e-13 PD=5.24e-06 PS=1.54e-06 $X=1390 $Y=2410 $dt=1
.ends NA2JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX1 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=4
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.44533e-13 AS=2.016e-13 PD=1.44667e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=6.6e-07 AD=2.88e-13 AS=3.84267e-13 PD=2.28e-06 PS=2.27333e-06 $X=1590 $Y=890 $dt=0
M2 vdd3i! A 6 vdd3i! pe3i L=3e-07 W=9e-07 AD=4.7931e-13 AS=4.32e-13 PD=1.95649e-06 PS=2.76e-06 $X=620 $Y=2410 $dt=1
M3 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=5.712e-13 AS=7.7739e-13 PD=3.70971e-06 PS=3.17322e-06 $X=1640 $Y=2410 $dt=1
.ends BUJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DFRRQJI3VX4                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DFRRQJI3VX4 vdd3i! gnd3i! RN D C Q
*.DEVICECLIMB
** N=23 EP=6 FDC=36
M0 gnd3i! 17 19 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=4.272e-13 PD=1.43e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 10 RN gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.28952e-13 AS=2.403e-13 PD=2.36956e-06 PS=1.43e-06 $X=1510 $Y=660 $dt=0
M2 18 19 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.55236e-13 PD=6.7e-07 PS=1.11822e-06 $X=2340 $Y=1390 $dt=0
M3 17 9 18 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=2940 $Y=1390 $dt=0
M4 16 15 17 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=3830 $Y=1390 $dt=0
M5 10 D 16 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.835e-13 AS=5.25e-14 PD=2.19e-06 PS=6.7e-07 $X=4430 $Y=1390 $dt=0
M6 gnd3i! C 15 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.659e-13 AS=2.016e-13 PD=1.21e-06 PS=1.8e-06 $X=6060 $Y=1390 $dt=0
M7 9 15 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.95e-13 AS=1.659e-13 PD=2.23e-06 PS=1.21e-06 $X=7045 $Y=1390 $dt=0
M8 14 19 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=8695 $Y=1020 $dt=0
M9 13 9 14 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=9295 $Y=1020 $dt=0
M10 12 15 13 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=10185 $Y=1020 $dt=0
M11 8 11 12 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.55817e-13 AS=5.25e-14 PD=9.68244e-07 PS=6.7e-07 $X=10785 $Y=1020 $dt=0
M12 gnd3i! RN 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.60325e-13 AS=3.30183e-13 PD=1.475e-06 PS=2.05176e-06 $X=11755 $Y=660 $dt=0
M13 11 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=2.60325e-13 PD=2.74e-06 PS=1.475e-06 $X=12690 $Y=660 $dt=0
M14 Q 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=4.272e-13 PD=1.43e-06 PS=2.74e-06 $X=14280 $Y=660 $dt=0
M15 gnd3i! 13 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=15170 $Y=660 $dt=0
M16 Q 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=16060 $Y=660 $dt=0
M17 gnd3i! 13 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=2.403e-13 PD=2.74e-06 PS=1.43e-06 $X=16950 $Y=660 $dt=0
M18 vdd3i! 17 19 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.54046e-13 AS=6.768e-13 PD=2.58169e-06 PS=3.78e-06 $X=620 $Y=2410 $dt=1
M19 17 RN vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.136e-13 AS=2.31854e-13 PD=2.4e-06 PS=1.31831e-06 $X=1460 $Y=2670 $dt=1
M20 23 19 vdd3i! vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=5.1875e-13 PD=6.7e-07 PS=2.99e-06 $X=3080 $Y=3400 $dt=1
M21 17 15 23 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=1.21617e-13 AS=5.25e-14 PD=9.13043e-07 PS=6.7e-07 $X=3630 $Y=3400 $dt=1
M22 22 9 17 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=1.2e-13 AS=2.77983e-13 PD=1.21e-06 PS=2.08696e-06 $X=4470 $Y=2860 $dt=1
M23 vdd3i! D 22 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=5.00229e-13 AS=1.2e-13 PD=2.34286e-06 PS=1.21e-06 $X=5020 $Y=2860 $dt=1
M24 15 C vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=4.94875e-13 AS=3.75171e-13 PD=3.04e-06 PS=1.75714e-06 $X=6060 $Y=2860 $dt=1
M25 vdd3i! 15 9 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.92547e-13 AS=3.528e-13 PD=1.8586e-06 PS=2.42e-06 $X=7720 $Y=2670 $dt=1
M26 21 19 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=1.25e-13 AS=5.45203e-13 PD=1.25e-06 PS=2.5814e-06 $X=8740 $Y=2820 $dt=1
M27 13 15 21 vdd3i! pe3i L=3e-07 W=1e-06 AD=2.96338e-13 AS=1.25e-13 PD=2.19718e-06 PS=1.25e-06 $X=9290 $Y=2820 $dt=1
M28 20 9 13 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=1.24462e-13 PD=6.7e-07 PS=9.22817e-07 $X=10150 $Y=3235 $dt=1
M29 vdd3i! 11 20 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=2.90656e-13 AS=5.25e-14 PD=1.25671e-06 PS=6.7e-07 $X=10700 $Y=3235 $dt=1
M30 vdd3i! RN 13 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=4.98268e-13 AS=2.976e-13 PD=2.15435e-06 PS=2.4e-06 $X=11900 $Y=2410 $dt=1
M31 11 13 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=9.75775e-13 PD=3.78e-06 PS=4.21894e-06 $X=12740 $Y=2410 $dt=1
M32 Q 13 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=1.1618e-12 PD=1.95e-06 PS=4.88e-06 $X=14480 $Y=2410 $dt=1
M33 vdd3i! 13 Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=3.807e-13 PD=1.95e-06 PS=1.95e-06 $X=15320 $Y=2410 $dt=1
M34 Q 13 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=3.807e-13 PD=1.95e-06 PS=1.95e-06 $X=16160 $Y=2410 $dt=1
M35 vdd3i! 13 Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=3.807e-13 PD=3.78e-06 PS=1.95e-06 $X=17000 $Y=2410 $dt=1
.ends DFRRQJI3VX4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX0                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX0 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=4
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.923e-13 AS=2.016e-13 PD=2.005e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=3.923e-13 PD=1.8e-06 PS=2.005e-06 $X=1735 $Y=1130 $dt=0
M2 vdd3i! A 6 vdd3i! pe3i L=3e-07 W=9e-07 AD=5.7805e-13 AS=4.32e-13 PD=2.33911e-06 PS=2.76e-06 $X=620 $Y=2410 $dt=1
M3 Q 6 vdd3i! vdd3i! pe3i L=3e-07 W=1.12e-06 AD=5.376e-13 AS=7.1935e-13 PD=3.2e-06 PS=2.91089e-06 $X=1785 $Y=2410 $dt=1
.ends BUJI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AN21JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AN21JI3VX1 vdd3i! gnd3i! B A Q C
*.DEVICECLIMB
** N=9 EP=6 FDC=6
M0 8 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=6.47e-13 PD=1.14e-06 PS=3.58e-06 $X=690 $Y=660 $dt=0
M1 Q A 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.28413e-13 AS=1.1125e-13 PD=1.78572e-06 PS=1.14e-06 $X=1290 $Y=660 $dt=0
M2 gnd3i! C Q gnd3i! ne3i L=3.5e-07 W=6.65e-07 AD=6.369e-13 AS=2.45387e-13 PD=3.6e-06 PS=1.33428e-06 $X=2310 $Y=885 $dt=0
M3 vdd3i! B 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.371e-13 AS=6.768e-13 PD=2.03e-06 PS=3.78e-06 $X=620 $Y=2410 $dt=1
M4 9 A vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=4.371e-13 PD=1.95e-06 PS=2.03e-06 $X=1540 $Y=2410 $dt=1
M5 Q C 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.614e-13 AS=3.807e-13 PD=3.9e-06 PS=1.95e-06 $X=2380 $Y=2410 $dt=1
.ends AN21JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: EN3JI3VX1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt EN3JI3VX1 vdd3i! gnd3i! C B A Q
*.DEVICECLIMB
** N=16 EP=6 FDC=20
M0 13 C gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=2.016e-13 PD=9.6e-07 PS=1.8e-06 $X=620 $Y=1030 $dt=0
M1 gnd3i! B 13 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.97668e-13 AS=1.134e-13 PD=1.24213e-06 PS=9.6e-07 $X=1510 $Y=1030 $dt=0
M2 12 C gnd3i! gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=6.5e-14 AS=2.44732e-13 PD=7.7e-07 PS=1.53787e-06 $X=2730 $Y=930 $dt=0
M3 11 B 12 gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=1.404e-13 AS=6.5e-14 PD=1.06e-06 PS=7.7e-07 $X=3330 $Y=930 $dt=0
M4 gnd3i! 13 11 gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=5.308e-13 AS=1.404e-13 PD=3.32e-06 PS=1.06e-06 $X=4220 $Y=930 $dt=0
M5 9 11 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=5850 $Y=970 $dt=0
M6 gnd3i! A 9 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=6450 $Y=970 $dt=0
M7 8 A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=1.134e-13 PD=9.6e-07 PS=9.6e-07 $X=7340 $Y=970 $dt=0
M8 gnd3i! 11 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.965e-13 AS=1.134e-13 PD=3.17071e-06 PS=9.6e-07 $X=8230 $Y=970 $dt=0
M9 Q 10 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=2.0035e-13 PD=1.8e-06 PS=1.77071e-06 $X=9670 $Y=1130 $dt=0
M10 16 C vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.115e-13 AS=7.1585e-13 PD=1.71e-06 PS=3.85e-06 $X=645 $Y=2410 $dt=1
M11 13 B 16 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=5.5365e-13 AS=2.115e-13 PD=3.83e-06 PS=1.71e-06 $X=1245 $Y=2410 $dt=1
M12 vdd3i! C 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.23e-13 AS=5.8645e-13 PD=2.01e-06 PS=3.83e-06 $X=2675 $Y=2410 $dt=1
M13 14 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=4.23e-13 PD=2e-06 PS=2.01e-06 $X=3575 $Y=2410 $dt=1
M14 11 13 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.1205e-13 AS=4.1595e-13 PD=3.83e-06 PS=2e-06 $X=4465 $Y=2410 $dt=1
M15 10 11 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=9.1545e-13 PD=2e-06 PS=4.61e-06 $X=6095 $Y=2410 $dt=1
M16 vdd3i! A 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.956e-13 AS=4.1595e-13 PD=2.63e-06 PS=2e-06 $X=6985 $Y=2410 $dt=1
M17 15 A vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.115e-13 AS=6.956e-13 PD=1.71e-06 PS=2.63e-06 $X=8155 $Y=2410 $dt=1
M18 Q 11 15 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.66787e-13 AS=2.115e-13 PD=2.36668e-06 PS=1.71e-06 $X=8755 $Y=2410 $dt=1
M19 vdd3i! 10 Q vdd3i! pe3i L=3e-07 W=9.85e-07 AD=8.62325e-13 AS=3.26088e-13 PD=4.61e-06 PS=1.65332e-06 $X=9655 $Y=2410 $dt=1
.ends EN3JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA3I2JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA3I2JI3VX1 vdd3i! gnd3i! AN BN C Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 9 AN gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=4.00432e-13 PD=9.6e-07 PS=2.10243e-06 $X=540 $Y=1130 $dt=0
M1 gnd3i! BN 9 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=4.00432e-13 AS=1.134e-13 PD=2.10243e-06 PS=9.6e-07 $X=1430 $Y=1130 $dt=0
M2 8 C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=8.48535e-13 PD=1.14e-06 PS=4.45514e-06 $X=2290 $Y=660 $dt=0
M3 Q 9 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.806e-13 AS=1.1125e-13 PD=2.86e-06 PS=1.14e-06 $X=2890 $Y=660 $dt=0
M4 10 AN 9 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=4.08e-13 PD=1.1e-06 PS=2.66e-06 $X=620 $Y=2410 $dt=1
M5 vdd3i! BN 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=7.38476e-13 AS=1.0625e-13 PD=3.31526e-06 PS=1.1e-06 $X=1170 $Y=2410 $dt=1
M6 vdd3i! C Q vdd3i! pe3i L=3.00037e-07 W=1.00071e-06 AD=8.69412e-13 AS=2.376e-13 PD=3.90308e-06 PS=1.49071e-06 $X=2170 $Y=2410 $dt=1
M7 Q 9 vdd3i! vdd3i! pe3i L=3.00037e-07 W=1.00071e-06 AD=2.376e-13 AS=8.69412e-13 PD=1.49071e-06 PS=3.90308e-06 $X=3010 $Y=2410 $dt=1
.ends NA3I2JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA22JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA22JI3VX1 vdd3i! gnd3i! A B C Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 9 A 10 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=2.688e-13 PD=8.1e-07 PS=2.08e-06 $X=620 $Y=990 $dt=0
M1 gnd3i! B 9 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=3.3376e-13 AS=7e-14 PD=1.56028e-06 PS=8.1e-07 $X=1220 $Y=990 $dt=0
M2 8 C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=5.3044e-13 PD=1.14e-06 PS=2.47972e-06 $X=2350 $Y=660 $dt=0
M3 Q 10 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=1.1125e-13 PD=2.74e-06 PS=1.14e-06 $X=2950 $Y=660 $dt=0
M4 10 A vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=7.66562e-13 PD=1.24e-06 PS=3.33273e-06 $X=510 $Y=2410 $dt=1
M5 vdd3i! B 10 vdd3i! pe3i L=3e-07 W=7e-07 AD=7.66562e-13 AS=1.89e-13 PD=3.33273e-06 PS=1.24e-06 $X=1350 $Y=2410 $dt=1
M6 vdd3i! C Q vdd3i! pe3i L=3.00052e-07 W=9.98995e-07 AD=1.09399e-12 AS=2.255e-13 PD=4.75626e-06 PS=1.46899e-06 $X=2190 $Y=2410 $dt=1
M7 Q 10 vdd3i! vdd3i! pe3i L=3.00052e-07 W=9.98995e-07 AD=2.255e-13 AS=1.09399e-12 PD=1.46899e-06 PS=4.75626e-06 $X=3030 $Y=2410 $dt=1
.ends NA22JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AN22JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AN22JI3VX1 vdd3i! gnd3i! B A Q C D
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 10 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=6.098e-13 PD=1.14e-06 PS=3.52e-06 $X=660 $Y=660 $dt=0
M1 Q A 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=1.1125e-13 PD=1.43e-06 PS=1.14e-06 $X=1260 $Y=660 $dt=0
M2 9 C Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=2.403e-13 PD=1.14e-06 PS=1.43e-06 $X=2150 $Y=660 $dt=0
M3 gnd3i! D 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=8.082e-13 AS=1.1125e-13 PD=3.84e-06 PS=1.14e-06 $X=2750 $Y=660 $dt=0
M4 vdd3i! B 11 vdd3i! pe3i L=3.01094e-07 W=1.47213e-06 AD=4.29e-13 AS=6.0945e-13 PD=2.32213e-06 PS=3.77213e-06 $X=660 $Y=2410 $dt=1
M5 11 A vdd3i! vdd3i! pe3i L=3.01094e-07 W=1.47213e-06 AD=4.05825e-13 AS=4.29e-13 PD=2.06213e-06 PS=2.32213e-06 $X=1310 $Y=2410 $dt=1
M6 Q C 11 vdd3i! pe3i L=3.01094e-07 W=1.47213e-06 AD=2.9925e-13 AS=4.05825e-13 PD=1.92213e-06 PS=2.06213e-06 $X=2200 $Y=2410 $dt=1
M7 11 D Q vdd3i! pe3i L=3.01094e-07 W=1.47213e-06 AD=6.252e-13 AS=2.9925e-13 PD=3.77213e-06 PS=1.92213e-06 $X=3100 $Y=2410 $dt=1
.ends AN22JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DLY1JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DLY1JI3VX1 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=8 EP=4 FDC=8
M0 gnd3i! A 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.591e-13 AS=2.016e-13 PD=2.13e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 6 8 gnd3i! gnd3i! ne3i L=8e-07 W=4.2e-07 AD=2.415e-13 AS=3.591e-13 PD=1.99e-06 PS=2.13e-06 $X=1590 $Y=1400 $dt=0
M2 gnd3i! 6 7 gnd3i! ne3i L=1e-06 W=4.2e-07 AD=2.6662e-13 AS=2.016e-13 PD=1.28565e-06 PS=1.8e-06 $X=2860 $Y=660 $dt=0
M3 Q 7 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.3165e-13 AS=5.6498e-13 PD=2.75e-06 PS=2.72435e-06 $X=4625 $Y=660 $dt=0
M4 vdd3i! A 8 vdd3i! pe3i L=3e-07 W=6.7e-07 AD=4.61962e-13 AS=3.3835e-13 PD=2.62468e-06 PS=2.35e-06 $X=645 $Y=2680 $dt=1
M5 6 8 vdd3i! vdd3i! pe3i L=1e-06 W=4.2e-07 AD=2.00088e-13 AS=2.89588e-13 PD=1.76778e-06 PS=1.64532e-06 $X=1590 $Y=2680 $dt=1
M6 vdd3i! 6 7 vdd3i! pe3i L=7.5e-07 W=4.2e-07 AD=2.78313e-13 AS=2.00088e-13 PD=1.17049e-06 PS=1.76778e-06 $X=3110 $Y=3400 $dt=1
M7 Q 7 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.191e-13 AS=9.34337e-13 PD=3.84e-06 PS=3.92951e-06 $X=4650 $Y=2410 $dt=1
.ends DLY1JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ON21JI3VX4                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ON21JI3VX4 vdd3i! gnd3i! B A C Q
*.DEVICECLIMB
** N=11 EP=6 FDC=16
M0 gnd3i! B 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=4.272e-13 PD=1.43e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 10 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=1510 $Y=660 $dt=0
M2 9 C 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.868e-13 AS=2.403e-13 PD=2.70971e-06 PS=1.43e-06 $X=2400 $Y=660 $dt=0
M3 gnd3i! 9 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.35783e-13 AS=4.34e-13 PD=1.42065e-06 PS=2.92971e-06 $X=3930 $Y=660 $dt=0
M4 Q 8 gnd3i! gnd3i! ne3i L=3.49164e-07 W=8.96213e-07 AD=2.32912e-13 AS=2.37429e-13 PD=1.42121e-06 PS=1.43057e-06 $X=4820 $Y=660 $dt=0
M5 gnd3i! 8 Q gnd3i! ne3i L=3.49164e-07 W=8.96213e-07 AD=2.32912e-13 AS=2.32912e-13 PD=1.42121e-06 PS=1.42121e-06 $X=5680 $Y=660 $dt=0
M6 Q 8 gnd3i! gnd3i! ne3i L=3.49164e-07 W=8.96213e-07 AD=2.32912e-13 AS=2.32912e-13 PD=1.42121e-06 PS=1.42121e-06 $X=6570 $Y=660 $dt=0
M7 gnd3i! 8 Q gnd3i! ne3i L=3.49164e-07 W=8.96213e-07 AD=4.19812e-13 AS=2.32912e-13 PD=2.73121e-06 PS=1.42121e-06 $X=7430 $Y=660 $dt=0
M8 11 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=9.418e-13 PD=1.66e-06 PS=4.63e-06 $X=695 $Y=2410 $dt=1
M9 9 A 11 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.68825e-13 AS=1.7625e-13 PD=2.075e-06 PS=1.66e-06 $X=1245 $Y=2410 $dt=1
M10 vdd3i! C 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.285e-12 AS=4.68825e-13 PD=5.02e-06 PS=2.075e-06 $X=2210 $Y=2410 $dt=1
M11 vdd3i! 9 8 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=5.48179e-13 AS=6.768e-13 PD=2.4141e-06 PS=3.78e-06 $X=4020 $Y=2410 $dt=1
M12 Q 8 vdd3i! vdd3i! pe3i L=3.00021e-07 W=1.42657e-06 AD=3.433e-13 AS=5.54621e-13 PD=1.92657e-06 PS=2.44247e-06 $X=4960 $Y=2410 $dt=1
M13 vdd3i! 8 Q vdd3i! pe3i L=3.00021e-07 W=1.42657e-06 AD=4.866e-13 AS=3.433e-13 PD=2.35657e-06 PS=1.92657e-06 $X=5800 $Y=2410 $dt=1
M14 Q 8 vdd3i! vdd3i! pe3i L=3.00021e-07 W=1.42657e-06 AD=3.433e-13 AS=4.866e-13 PD=1.92657e-06 PS=2.35657e-06 $X=6640 $Y=2410 $dt=1
M15 vdd3i! 8 Q vdd3i! pe3i L=3.00021e-07 W=1.42657e-06 AD=8.562e-13 AS=3.433e-13 PD=4.53657e-06 PS=1.92657e-06 $X=7480 $Y=2410 $dt=1
.ends ON21JI3VX4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INJI3VX6                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INJI3VX6 vdd3i! gnd3i! Q A
*.DEVICECLIMB
** N=5 EP=4 FDC=10
M0 gnd3i! A Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=4.272e-13 PD=1.86e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=1590 $Y=660 $dt=0
M2 gnd3i! A Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.114e-13 AS=2.403e-13 PD=1.96e-06 PS=1.43e-06 $X=2480 $Y=660 $dt=0
M3 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=4.114e-13 PD=2.74e-06 PS=1.96e-06 $X=3550 $Y=660 $dt=0
M4 Q A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=5.79287e-13 PD=1.86506e-06 PS=3.69506e-06 $X=475 $Y=2410 $dt=1
M5 vdd3i! A Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1315 $Y=2410 $dt=1
M6 Q A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1865 $Y=2410 $dt=1
M7 vdd3i! A Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=2705 $Y=2410 $dt=1
M8 Q A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=3255 $Y=2410 $dt=1
M9 vdd3i! A Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=1.01149e-12 AS=2.54913e-13 PD=4.73506e-06 PS=1.86506e-06 $X=4095 $Y=2410 $dt=1
.ends INJI3VX6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA3I1JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA3I1JI3VX1 vdd3i! gnd3i! AN Q B C
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 gnd3i! AN 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.40779e-13 AS=2.016e-13 PD=1.24397e-06 PS=1.8e-06 $X=620 $Y=660 $dt=0
M1 9 10 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.26825e-13 AS=5.10221e-13 PD=1.175e-06 PS=2.63603e-06 $X=1670 $Y=660 $dt=0
M2 8 B 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.31275e-13 AS=1.26825e-13 PD=1.185e-06 PS=1.175e-06 $X=2305 $Y=660 $dt=0
M3 Q C 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=1.31275e-13 PD=2.74e-06 PS=1.185e-06 $X=2950 $Y=660 $dt=0
M4 vdd3i! AN 10 vdd3i! pe3i L=3e-07 W=7e-07 AD=4.82246e-13 AS=3.36e-13 PD=2.26063e-06 PS=2.36e-06 $X=620 $Y=2410 $dt=1
M5 vdd3i! 10 Q vdd3i! pe3i L=3.00059e-07 W=1.00314e-06 AD=6.91085e-13 AS=2.195e-13 PD=3.2396e-06 PS=1.46314e-06 $X=1430 $Y=2410 $dt=1
M6 Q B vdd3i! vdd3i! pe3i L=3.00059e-07 W=1.00314e-06 AD=2.195e-13 AS=6.91085e-13 PD=1.46314e-06 PS=3.2396e-06 $X=2270 $Y=2410 $dt=1
M7 Q C vdd3i! vdd3i! pe3i L=3.00059e-07 W=1.00314e-06 AD=4.232e-13 AS=6.91085e-13 PD=2.85314e-06 PS=3.2396e-06 $X=3000 $Y=2410 $dt=1
.ends NA3I1JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX8                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX8 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=19
M0 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=6.098e-13 PD=1.43e-06 PS=3.52e-06 $X=660 $Y=660 $dt=0
M1 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.804e-13 AS=2.403e-13 PD=1.91e-06 PS=1.43e-06 $X=1550 $Y=660 $dt=0
M2 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.804e-13 PD=1.43e-06 PS=1.91e-06 $X=2570 $Y=660 $dt=0
M3 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=3460 $Y=660 $dt=0
M4 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=4430 $Y=660 $dt=0
M5 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=5320 $Y=660 $dt=0
M6 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=6290 $Y=660 $dt=0
M7 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=8.702e-13 AS=2.403e-13 PD=3.94e-06 PS=1.43e-06 $X=7180 $Y=660 $dt=0
M8 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=5.51013e-13 PD=1.86506e-06 PS=3.69506e-06 $X=620 $Y=2410 $dt=1
M9 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.61963e-13 AS=2.83187e-13 PD=1.87506e-06 PS=1.86506e-06 $X=1170 $Y=2410 $dt=1
M10 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.61963e-13 PD=1.86506e-06 PS=1.87506e-06 $X=2020 $Y=2410 $dt=1
M11 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.61963e-13 AS=2.83187e-13 PD=1.87506e-06 PS=1.86506e-06 $X=2570 $Y=2410 $dt=1
M12 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.61963e-13 PD=1.86506e-06 PS=1.87506e-06 $X=3420 $Y=2410 $dt=1
M13 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.61963e-13 AS=2.83187e-13 PD=1.87506e-06 PS=1.86506e-06 $X=3970 $Y=2410 $dt=1
M14 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.61963e-13 PD=1.86506e-06 PS=1.87506e-06 $X=4820 $Y=2410 $dt=1
M15 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.61963e-13 AS=2.83187e-13 PD=1.87506e-06 PS=1.86506e-06 $X=5370 $Y=2410 $dt=1
M16 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.61963e-13 PD=1.86506e-06 PS=1.87506e-06 $X=6220 $Y=2410 $dt=1
M17 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.61963e-13 AS=2.83187e-13 PD=1.87506e-06 PS=1.86506e-06 $X=6770 $Y=2410 $dt=1
M18 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=5.79287e-13 AS=2.61963e-13 PD=3.69506e-06 PS=1.87506e-06 $X=7620 $Y=2410 $dt=1
.ends BUJI3VX8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DFRRQJI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DFRRQJI3VX1 vdd3i! gnd3i! RN D C Q
*.DEVICECLIMB
** N=23 EP=6 FDC=30
M0 gnd3i! 17 19 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.39017e-13 AS=2.016e-13 PD=9.16947e-07 PS=1.8e-06 $X=620 $Y=660 $dt=0
M1 10 RN gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.28952e-13 AS=2.94583e-13 PD=2.36956e-06 PS=1.94305e-06 $X=1510 $Y=660 $dt=0
M2 18 19 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.55236e-13 PD=6.7e-07 PS=1.11822e-06 $X=2340 $Y=1390 $dt=0
M3 17 9 18 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=2940 $Y=1390 $dt=0
M4 16 15 17 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=3830 $Y=1390 $dt=0
M5 10 D 16 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.835e-13 AS=5.25e-14 PD=2.19e-06 PS=6.7e-07 $X=4430 $Y=1390 $dt=0
M6 gnd3i! C 15 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.659e-13 AS=2.016e-13 PD=1.21e-06 PS=1.8e-06 $X=6060 $Y=1390 $dt=0
M7 9 15 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.95e-13 AS=1.659e-13 PD=2.23e-06 PS=1.21e-06 $X=7045 $Y=1390 $dt=0
M8 14 19 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=8695 $Y=1020 $dt=0
M9 13 9 14 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=9295 $Y=1020 $dt=0
M10 12 15 13 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=10185 $Y=1020 $dt=0
M11 8 11 12 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.55817e-13 AS=5.25e-14 PD=9.68244e-07 PS=6.7e-07 $X=10785 $Y=1020 $dt=0
M12 gnd3i! RN 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=6.52289e-13 AS=3.30183e-13 PD=3.3375e-06 PS=2.05176e-06 $X=11755 $Y=660 $dt=0
M13 11 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=3.07822e-13 PD=1.8e-06 PS=1.575e-06 $X=12560 $Y=1130 $dt=0
M14 Q 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=6.52289e-13 PD=2.74e-06 PS=3.3375e-06 $X=14150 $Y=660 $dt=0
M15 vdd3i! 17 19 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=1.944e-13 AS=3.456e-13 PD=1.26e-06 PS=2.4e-06 $X=620 $Y=2670 $dt=1
M16 17 RN vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.136e-13 AS=1.944e-13 PD=2.4e-06 PS=1.26e-06 $X=1460 $Y=2670 $dt=1
M17 23 19 vdd3i! vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=5.1875e-13 PD=6.7e-07 PS=2.99e-06 $X=3080 $Y=3400 $dt=1
M18 17 15 23 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=1.21617e-13 AS=5.25e-14 PD=9.13043e-07 PS=6.7e-07 $X=3630 $Y=3400 $dt=1
M19 22 9 17 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=1.2e-13 AS=2.77983e-13 PD=1.21e-06 PS=2.08696e-06 $X=4470 $Y=2860 $dt=1
M20 vdd3i! D 22 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=5.00229e-13 AS=1.2e-13 PD=2.34286e-06 PS=1.21e-06 $X=5020 $Y=2860 $dt=1
M21 15 C vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=4.94875e-13 AS=3.75171e-13 PD=3.04e-06 PS=1.75714e-06 $X=6060 $Y=2860 $dt=1
M22 vdd3i! 15 9 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.92547e-13 AS=3.528e-13 PD=1.8586e-06 PS=2.42e-06 $X=7720 $Y=2670 $dt=1
M23 21 19 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=1.25e-13 AS=5.45203e-13 PD=1.25e-06 PS=2.5814e-06 $X=8740 $Y=2820 $dt=1
M24 13 15 21 vdd3i! pe3i L=3e-07 W=1e-06 AD=2.96338e-13 AS=1.25e-13 PD=2.19718e-06 PS=1.25e-06 $X=9290 $Y=2820 $dt=1
M25 20 9 13 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=1.24462e-13 PD=6.7e-07 PS=9.22817e-07 $X=10150 $Y=3235 $dt=1
M26 vdd3i! 11 20 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=4.10996e-13 AS=5.25e-14 PD=1.64789e-06 PS=6.7e-07 $X=10700 $Y=3235 $dt=1
M27 vdd3i! RN 13 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=7.04565e-13 AS=2.976e-13 PD=2.82495e-06 PS=2.4e-06 $X=11900 $Y=2410 $dt=1
M28 11 13 vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.456e-13 AS=7.04565e-13 PD=2.4e-06 PS=2.82495e-06 $X=12740 $Y=2410 $dt=1
M29 Q 13 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=1.37977e-12 PD=3.78e-06 PS=5.5322e-06 $X=14200 $Y=2410 $dt=1
.ends DFRRQJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ON211JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ON211JI3VX1 vdd3i! gnd3i! B Q A C D
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 Q B 10 gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.27987e-13 AS=4.20337e-13 PD=1.41536e-06 PS=2.75536e-06 $X=620 $Y=660 $dt=0
M1 10 A Q gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.30287e-13 AS=2.27987e-13 PD=1.43036e-06 PS=1.41536e-06 $X=1460 $Y=660 $dt=0
M2 9 C 10 gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=1.21188e-13 AS=2.30287e-13 PD=1.17536e-06 PS=1.43036e-06 $X=2350 $Y=660 $dt=0
M3 gnd3i! D 9 gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=4.20337e-13 AS=1.21188e-13 PD=2.75536e-06 PS=1.17536e-06 $X=2950 $Y=660 $dt=0
M4 11 B vdd3i! vdd3i! pe3i L=3e-07 W=1.38e-06 AD=1.725e-13 AS=9.388e-13 PD=1.63e-06 PS=4.63e-06 $X=695 $Y=2410 $dt=1
M5 Q A 11 vdd3i! pe3i L=3e-07 W=1.38e-06 AD=4.69617e-13 AS=1.725e-13 PD=2.38255e-06 PS=1.63e-06 $X=1245 $Y=2410 $dt=1
M6 vdd3i! C Q vdd3i! pe3i L=3.00049e-07 W=9.66924e-07 AD=4.25413e-13 AS=3.29046e-13 PD=2.34192e-06 PS=1.66938e-06 $X=2210 $Y=2410 $dt=1
M7 Q D vdd3i! vdd3i! pe3i L=3.00049e-07 W=9.66924e-07 AD=4.20162e-13 AS=4.25413e-13 PD=2.80192e-06 PS=2.34192e-06 $X=3000 $Y=2410 $dt=1
.ends ON211JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ON22JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ON22JI3VX1 vdd3i! gnd3i! D C Q A B
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 gnd3i! D 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=4.272e-13 PD=1.86e-06 PS=2.74e-06 $X=720 $Y=660 $dt=0
M1 9 C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=1690 $Y=660 $dt=0
M2 Q A 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=2580 $Y=660 $dt=0
M3 9 B Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.666e-13 AS=2.403e-13 PD=2.84e-06 PS=1.43e-06 $X=3470 $Y=660 $dt=0
M4 11 D vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=8.802e-13 PD=1.66e-06 PS=4.56e-06 $X=1120 $Y=2410 $dt=1
M5 Q C 11 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=1.7625e-13 PD=1.95e-06 PS=1.66e-06 $X=1670 $Y=2410 $dt=1
M6 10 A Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=3.807e-13 PD=1.66e-06 PS=1.95e-06 $X=2510 $Y=2410 $dt=1
M7 vdd3i! B 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=8.802e-13 AS=1.7625e-13 PD=4.56e-06 PS=1.66e-06 $X=3060 $Y=2410 $dt=1
.ends ON22JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DFRRQJI3VX2                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DFRRQJI3VX2 vdd3i! gnd3i! RN D C Q
*.DEVICECLIMB
** N=23 EP=6 FDC=32
M0 gnd3i! 17 19 gnd3i! ne3i L=3.5e-07 W=6.6e-07 AD=1.94849e-13 AS=3.168e-13 PD=1.21781e-06 PS=2.28e-06 $X=620 $Y=660 $dt=0
M1 10 RN gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.28952e-13 AS=2.62751e-13 PD=2.36956e-06 PS=1.64219e-06 $X=1510 $Y=660 $dt=0
M2 18 19 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.55236e-13 PD=6.7e-07 PS=1.11822e-06 $X=2340 $Y=1390 $dt=0
M3 17 9 18 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=2940 $Y=1390 $dt=0
M4 16 15 17 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=3830 $Y=1390 $dt=0
M5 10 D 16 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.835e-13 AS=5.25e-14 PD=2.19e-06 PS=6.7e-07 $X=4430 $Y=1390 $dt=0
M6 gnd3i! C 15 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.659e-13 AS=2.016e-13 PD=1.21e-06 PS=1.8e-06 $X=6060 $Y=1390 $dt=0
M7 9 15 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.95e-13 AS=1.659e-13 PD=2.23e-06 PS=1.21e-06 $X=7045 $Y=1390 $dt=0
M8 14 19 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=8695 $Y=1020 $dt=0
M9 13 9 14 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=9295 $Y=1020 $dt=0
M10 12 15 13 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=10185 $Y=1020 $dt=0
M11 8 11 12 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.55817e-13 AS=5.25e-14 PD=9.68244e-07 PS=6.7e-07 $X=10785 $Y=1020 $dt=0
M12 gnd3i! RN 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=5.94987e-13 AS=3.30183e-13 PD=3.35209e-06 PS=2.05176e-06 $X=11755 $Y=660 $dt=0
M13 11 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=6.6e-07 AD=3.168e-13 AS=4.41226e-13 PD=2.28e-06 PS=2.48582e-06 $X=12750 $Y=890 $dt=0
M14 Q 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=5.94987e-13 PD=1.43e-06 PS=3.35209e-06 $X=14380 $Y=660 $dt=0
M15 gnd3i! 13 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=2.403e-13 PD=2.74e-06 PS=1.43e-06 $X=15270 $Y=660 $dt=0
M16 vdd3i! 17 19 vdd3i! pe3i L=3e-07 W=1e-06 AD=2.97674e-13 AS=4.8e-13 PD=1.7907e-06 PS=2.96e-06 $X=620 $Y=2670 $dt=1
M17 17 RN vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.136e-13 AS=2.14326e-13 PD=2.4e-06 PS=1.2893e-06 $X=1460 $Y=2670 $dt=1
M18 23 19 vdd3i! vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=5.1875e-13 PD=6.7e-07 PS=2.99e-06 $X=3080 $Y=3400 $dt=1
M19 17 15 23 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=1.21617e-13 AS=5.25e-14 PD=9.13043e-07 PS=6.7e-07 $X=3630 $Y=3400 $dt=1
M20 22 9 17 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=1.2e-13 AS=2.77983e-13 PD=1.21e-06 PS=2.08696e-06 $X=4470 $Y=2860 $dt=1
M21 vdd3i! D 22 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=5.00229e-13 AS=1.2e-13 PD=2.34286e-06 PS=1.21e-06 $X=5020 $Y=2860 $dt=1
M22 15 C vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=4.56625e-13 AS=3.75171e-13 PD=2.86e-06 PS=1.75714e-06 $X=6060 $Y=2860 $dt=1
M23 vdd3i! 15 9 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.92547e-13 AS=3.528e-13 PD=1.8586e-06 PS=2.42e-06 $X=7720 $Y=2670 $dt=1
M24 21 19 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=1.25e-13 AS=5.45203e-13 PD=1.25e-06 PS=2.5814e-06 $X=8740 $Y=2820 $dt=1
M25 13 15 21 vdd3i! pe3i L=3e-07 W=1e-06 AD=2.96338e-13 AS=1.25e-13 PD=2.19718e-06 PS=1.25e-06 $X=9290 $Y=2820 $dt=1
M26 20 9 13 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=1.24462e-13 PD=6.7e-07 PS=9.22817e-07 $X=10150 $Y=3235 $dt=1
M27 vdd3i! 11 20 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=3.93439e-13 AS=5.25e-14 PD=1.64096e-06 PS=6.7e-07 $X=10700 $Y=3235 $dt=1
M28 vdd3i! RN 13 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=6.74468e-13 AS=2.976e-13 PD=2.81307e-06 PS=2.4e-06 $X=11900 $Y=2410 $dt=1
M29 11 13 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=4.8e-13 AS=9.36761e-13 PD=2.96e-06 PS=3.90704e-06 $X=12740 $Y=2410 $dt=1
M30 Q 13 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=1.32083e-12 PD=1.95e-06 PS=5.50893e-06 $X=14440 $Y=2410 $dt=1
M31 vdd3i! 13 Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=8.802e-13 AS=3.807e-13 PD=4.56e-06 PS=1.95e-06 $X=15280 $Y=2410 $dt=1
.ends DFRRQJI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: EO3JI3VX1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt EO3JI3VX1 vdd3i! gnd3i! C B A Q
*.DEVICECLIMB
** N=16 EP=6 FDC=20
M0 12 C gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.628e-13 PD=9.6e-07 PS=3.52e-06 $X=660 $Y=1130 $dt=0
M1 gnd3i! B 12 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.30196e-13 AS=1.134e-13 PD=1.36723e-06 PS=9.6e-07 $X=1550 $Y=1130 $dt=0
M2 11 C gnd3i! gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=6.5e-14 AS=2.85004e-13 PD=7.7e-07 PS=1.69277e-06 $X=2910 $Y=1030 $dt=0
M3 10 B 11 gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=1.404e-13 AS=6.5e-14 PD=1.06e-06 PS=7.7e-07 $X=3510 $Y=1030 $dt=0
M4 gnd3i! 12 10 gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=8.05779e-13 AS=1.404e-13 PD=2.83787e-06 PS=1.06e-06 $X=4400 $Y=1030 $dt=0
M5 9 10 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=6.50821e-13 PD=9.6e-07 PS=2.29213e-06 $X=6075 $Y=1130 $dt=0
M6 gnd3i! A 9 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.90537e-13 AS=1.134e-13 PD=1.53255e-06 PS=9.6e-07 $X=6965 $Y=1130 $dt=0
M7 8 A gnd3i! gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=6.5e-14 AS=3.59713e-13 PD=7.7e-07 PS=1.89745e-06 $X=8140 $Y=1030 $dt=0
M8 Q 10 8 gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=1.404e-13 AS=6.5e-14 PD=1.06e-06 PS=7.7e-07 $X=8740 $Y=1030 $dt=0
M9 gnd3i! 9 Q gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=5.728e-13 AS=1.404e-13 PD=3.52e-06 PS=1.06e-06 $X=9630 $Y=1030 $dt=0
M10 16 C vdd3i! vdd3i! pe3i L=3e-07 W=1.3e-06 AD=1.95e-13 AS=6.603e-13 PD=1.6e-06 PS=3.63e-06 $X=645 $Y=2520 $dt=1
M11 12 B 16 vdd3i! pe3i L=3e-07 W=1.3e-06 AD=5.157e-13 AS=1.95e-13 PD=3.61e-06 PS=1.6e-06 $X=1245 $Y=2520 $dt=1
M12 vdd3i! C 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=5.8645e-13 PD=2e-06 PS=3.83e-06 $X=2675 $Y=2410 $dt=1
M13 14 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=4.1595e-13 PD=2e-06 PS=2e-06 $X=3565 $Y=2410 $dt=1
M14 10 12 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=5.6965e-13 AS=4.1595e-13 PD=3.83e-06 PS=2e-06 $X=4455 $Y=2410 $dt=1
M15 15 10 vdd3i! vdd3i! pe3i L=3e-07 W=1.3e-06 AD=1.95e-13 AS=5.301e-13 PD=1.6e-06 PS=3.61e-06 $X=5885 $Y=2410 $dt=1
M16 9 A 15 vdd3i! pe3i L=3e-07 W=1.3e-06 AD=5.157e-13 AS=1.95e-13 PD=3.61e-06 PS=1.6e-06 $X=6485 $Y=2410 $dt=1
M17 vdd3i! A 13 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=5.8645e-13 PD=2e-06 PS=3.83e-06 $X=7915 $Y=2410 $dt=1
M18 13 10 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=4.1595e-13 PD=2e-06 PS=2e-06 $X=8805 $Y=2410 $dt=1
M19 Q 9 13 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.1205e-13 AS=4.1595e-13 PD=3.83e-06 PS=2e-06 $X=9695 $Y=2410 $dt=1
.ends EO3JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO2JI3VX0 vdd3i! gnd3i! B Q A
*.DEVICECLIMB
** N=7 EP=5 FDC=4
M0 Q B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=7.244e-13 PD=9.6e-07 PS=4.14e-06 $X=500 $Y=1130 $dt=0
M1 gnd3i! A Q gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=7.244e-13 AS=1.134e-13 PD=4.14e-06 PS=9.6e-07 $X=1390 $Y=1130 $dt=0
M2 7 B vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=9.298e-13 PD=1.1e-06 PS=4.68e-06 $X=720 $Y=2410 $dt=1
M3 Q A 7 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.08e-13 AS=1.0625e-13 PD=2.66e-06 PS=1.1e-06 $X=1270 $Y=2410 $dt=1
.ends NO2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ON21JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ON21JI3VX1 vdd3i! gnd3i! B A Q C
*.DEVICECLIMB
** N=9 EP=6 FDC=6
M0 gnd3i! B 8 gnd3i! ne3i L=3.4958e-07 W=8.92071e-07 AD=2.40125e-13 AS=4.24712e-13 PD=1.43207e-06 PS=2.73707e-06 $X=615 $Y=660 $dt=0
M1 8 A gnd3i! gnd3i! ne3i L=3.4958e-07 W=8.92071e-07 AD=2.37987e-13 AS=2.40125e-13 PD=1.42707e-06 PS=1.43207e-06 $X=1505 $Y=660 $dt=0
M2 Q C 8 gnd3i! ne3i L=3.4958e-07 W=8.92071e-07 AD=4.24712e-13 AS=2.37987e-13 PD=2.73707e-06 PS=1.42707e-06 $X=2395 $Y=660 $dt=0
M3 9 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=9.418e-13 PD=1.66e-06 PS=4.63e-06 $X=695 $Y=2410 $dt=1
M4 Q A 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.75706e-13 AS=1.7625e-13 PD=2.44322e-06 PS=1.66e-06 $X=1245 $Y=2410 $dt=1
M5 vdd3i! C Q vdd3i! pe3i L=3e-07 W=9.85e-07 AD=1.1721e-12 AS=3.32319e-13 PD=4.94e-06 PS=1.70678e-06 $X=2210 $Y=2410 $dt=1
.ends ON21JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OR4JI3VX1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OR4JI3VX1 vdd3i! gnd3i! C D Q B A
*.DEVICECLIMB
** N=13 EP=7 FDC=12
M0 11 C gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=4.12474e-13 PD=9.6e-07 PS=2.12185e-06 $X=510 $Y=1130 $dt=0
M1 gnd3i! D 11 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=4.12474e-13 AS=1.134e-13 PD=2.12185e-06 PS=9.6e-07 $X=1400 $Y=1130 $dt=0
M2 10 11 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=8.74052e-13 PD=1.14e-06 PS=4.4963e-06 $X=2330 $Y=660 $dt=0
M3 Q 9 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.56e-13 AS=1.1125e-13 PD=2.64627e-06 PS=1.14e-06 $X=2930 $Y=660 $dt=0
M4 9 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=7.908e-13 PD=9.6e-07 PS=4.27314e-06 $X=4410 $Y=1130 $dt=0
M5 gnd3i! A 9 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=7.908e-13 AS=1.134e-13 PD=4.27314e-06 PS=9.6e-07 $X=5300 $Y=1130 $dt=0
M6 13 C 11 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=4.08e-13 PD=1.1e-06 PS=2.66e-06 $X=620 $Y=2410 $dt=1
M7 vdd3i! D 13 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=6.21177e-13 AS=1.0625e-13 PD=2.08363e-06 PS=1.1e-06 $X=1170 $Y=2410 $dt=1
M8 Q 11 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=1.03042e-12 PD=1.95e-06 PS=3.45637e-06 $X=2480 $Y=2410 $dt=1
M9 vdd3i! 9 Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.09631e-12 AS=3.807e-13 PD=3.53124e-06 PS=1.95e-06 $X=3320 $Y=2410 $dt=1
M10 12 B vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=6.60894e-13 PD=1.1e-06 PS=2.12876e-06 $X=4690 $Y=2410 $dt=1
M11 9 A 12 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.08e-13 AS=1.0625e-13 PD=2.66e-06 PS=1.1e-06 $X=5240 $Y=2410 $dt=1
.ends OR4JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX16                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX16 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=39
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=4.272e-13 PD=1.43e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=1510 $Y=660 $dt=0
M2 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=2400 $Y=660 $dt=0
M3 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=3290 $Y=660 $dt=0
M4 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=4180 $Y=660 $dt=0
M5 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.4475e-13 AS=2.403e-13 PD=1.44e-06 PS=1.43e-06 $X=5070 $Y=660 $dt=0
M6 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.63267e-13 AS=2.4475e-13 PD=1.95905e-06 PS=1.44e-06 $X=5970 $Y=660 $dt=0
M7 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.26533e-13 PD=1.34e-06 PS=1.76095e-06 $X=6940 $Y=750 $dt=0
M8 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=7830 $Y=750 $dt=0
M9 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=8800 $Y=750 $dt=0
M10 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=9690 $Y=750 $dt=0
M11 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=10660 $Y=750 $dt=0
M12 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=11550 $Y=750 $dt=0
M13 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=12520 $Y=750 $dt=0
M14 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=13410 $Y=750 $dt=0
M15 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=14380 $Y=750 $dt=0
M16 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.84e-13 AS=2.16e-13 PD=2.56e-06 PS=1.34e-06 $X=15270 $Y=750 $dt=0
M17 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=5.79287e-13 PD=1.86506e-06 PS=3.69506e-06 $X=475 $Y=2410 $dt=1
M18 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1315 $Y=2410 $dt=1
M19 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1865 $Y=2410 $dt=1
M20 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=2705 $Y=2410 $dt=1
M21 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=3255 $Y=2410 $dt=1
M22 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=4095 $Y=2410 $dt=1
M23 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=4645 $Y=2410 $dt=1
M24 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=5485 $Y=2410 $dt=1
M25 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=6035 $Y=2410 $dt=1
M26 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=6875 $Y=2410 $dt=1
M27 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=7425 $Y=2410 $dt=1
M28 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=8265 $Y=2410 $dt=1
M29 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=8815 $Y=2410 $dt=1
M30 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=9655 $Y=2410 $dt=1
M31 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=10205 $Y=2410 $dt=1
M32 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=11045 $Y=2410 $dt=1
M33 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=11595 $Y=2410 $dt=1
M34 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=12435 $Y=2410 $dt=1
M35 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=12985 $Y=2410 $dt=1
M36 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=13825 $Y=2410 $dt=1
M37 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=14375 $Y=2410 $dt=1
M38 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=1.15229e-12 AS=2.54913e-13 PD=4.89506e-06 PS=1.86506e-06 $X=15215 $Y=2410 $dt=1
.ends BUJI3VX16

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX6                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX6 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=14
M0 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=6.008e-13 PD=1.34e-06 PS=3.52e-06 $X=660 $Y=750 $dt=0
M1 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=5.84805e-13 AS=2.16e-13 PD=2.17751e-06 PS=1.34e-06 $X=1550 $Y=750 $dt=0
M2 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=6.50595e-13 PD=1.43e-06 PS=2.42249e-06 $X=2960 $Y=660 $dt=0
M3 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=3850 $Y=660 $dt=0
M4 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=4820 $Y=660 $dt=0
M5 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=6.098e-13 AS=2.403e-13 PD=3.52e-06 PS=1.43e-06 $X=5710 $Y=660 $dt=0
M6 6 A vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=6.3285e-13 PD=1.87971e-06 PS=3.75971e-06 $X=525 $Y=2410 $dt=1
M7 vdd3i! A 6 vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=3.7905e-13 AS=2.751e-13 PD=1.98971e-06 PS=1.87971e-06 $X=1365 $Y=2410 $dt=1
M8 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=3.7905e-13 PD=1.87971e-06 PS=1.98971e-06 $X=2075 $Y=2410 $dt=1
M9 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=3.3675e-13 AS=2.751e-13 PD=1.92971e-06 PS=1.87971e-06 $X=2915 $Y=2410 $dt=1
M10 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=3.3675e-13 PD=1.87971e-06 PS=1.92971e-06 $X=3565 $Y=2410 $dt=1
M11 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=3.3675e-13 AS=2.751e-13 PD=1.92971e-06 PS=1.87971e-06 $X=4405 $Y=2410 $dt=1
M12 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=3.3675e-13 PD=1.87971e-06 PS=1.92971e-06 $X=5055 $Y=2410 $dt=1
M13 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=6.3285e-13 AS=2.751e-13 PD=3.75971e-06 PS=1.87971e-06 $X=5895 $Y=2410 $dt=1
.ends BUJI3VX6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ON31JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ON31JI3VX1 vdd3i! gnd3i! A B C Q D
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 9 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=6.098e-13 PD=1.43e-06 PS=3.52e-06 $X=660 $Y=660 $dt=0
M1 gnd3i! B 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=1550 $Y=660 $dt=0
M2 9 C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=2520 $Y=660 $dt=0
M3 Q D 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=2.403e-13 PD=2.74e-06 PS=1.43e-06 $X=3410 $Y=660 $dt=0
M4 11 A vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=9.066e-13 PD=1.72e-06 PS=4.59e-06 $X=1145 $Y=2410 $dt=1
M5 10 B 11 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=2.1855e-13 PD=1.72e-06 PS=1.72e-06 $X=1755 $Y=2410 $dt=1
M6 Q C 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=5.30442e-13 AS=2.1855e-13 PD=2.60067e-06 PS=1.72e-06 $X=2365 $Y=2410 $dt=1
M7 vdd3i! D Q vdd3i! pe3i L=3e-07 W=8.4e-07 AD=1.1576e-12 AS=3.16008e-13 PD=4.94e-06 PS=1.54933e-06 $X=3330 $Y=2410 $dt=1
.ends ON31JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DLY4JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DLY4JI3VX1 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=12 EP=4 FDC=12
M0 gnd3i! A 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.323e-13 AS=2.016e-13 PD=1.05e-06 PS=1.8e-06 $X=620 $Y=660 $dt=0
M1 8 10 gnd3i! gnd3i! ne3i L=1.8e-06 W=4.2e-07 AD=1.736e-13 AS=1.323e-13 PD=1.58e-06 PS=1.05e-06 $X=1600 $Y=660 $dt=0
M2 8 10 9 gnd3i! ne3i L=1.8e-06 W=4.2e-07 AD=1.736e-13 AS=2.00088e-13 PD=1.58e-06 PS=1.76778e-06 $X=1600 $Y=1360 $dt=0
M3 gnd3i! 9 7 gnd3i! ne3i L=1.1e-06 W=4.2e-07 AD=4.30324e-13 AS=2.16e-13 PD=1.75053e-06 PS=1.66e-06 $X=4630 $Y=660 $dt=0
M4 6 9 7 gnd3i! ne3i L=1.1e-06 W=4.2e-07 AD=2.00088e-13 AS=2.16e-13 PD=1.76778e-06 PS=1.66e-06 $X=4630 $Y=1400 $dt=0
M5 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.4055e-13 AS=9.11876e-13 PD=2.77e-06 PS=3.70947e-06 $X=7220 $Y=660 $dt=0
M6 vdd3i! A 10 vdd3i! pe3i L=3e-07 W=7e-07 AD=5.26875e-13 AS=3.535e-13 PD=3.30625e-06 PS=2.41e-06 $X=645 $Y=2680 $dt=1
M7 12 10 9 vdd3i! pe3i L=1.2e-06 W=4.2e-07 AD=1.674e-13 AS=2.016e-13 PD=1.56e-06 PS=1.8e-06 $X=2100 $Y=2680 $dt=1
M8 12 10 vdd3i! vdd3i! pe3i L=1.2e-06 W=4.2e-07 AD=1.674e-13 AS=3.16125e-13 PD=1.56e-06 PS=1.98375e-06 $X=2100 $Y=3400 $dt=1
M9 6 9 11 vdd3i! pe3i L=1.9e-06 W=4.2e-07 AD=2.016e-13 AS=1.674e-13 PD=1.8e-06 PS=1.56e-06 $X=4220 $Y=2680 $dt=1
M10 vdd3i! 9 11 vdd3i! pe3i L=1.9e-06 W=4.2e-07 AD=2.6367e-13 AS=1.674e-13 PD=1.32426e-06 PS=1.56e-06 $X=4220 $Y=3400 $dt=1
M11 Q 6 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.332e-13 AS=8.8518e-13 PD=3.86e-06 PS=4.44574e-06 $X=7245 $Y=2410 $dt=1
.ends DLY4JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO2I1JI3VX2                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO2I1JI3VX2 vdd3i! gnd3i! AN Q B
*.DEVICECLIMB
** N=9 EP=5 FDC=10
M0 gnd3i! AN 7 gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.3695e-13 AS=4.15012e-13 PD=1.44536e-06 PS=2.72536e-06 $X=595 $Y=660 $dt=0
M1 Q 7 gnd3i! gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.28113e-13 AS=2.3695e-13 PD=1.41536e-06 PS=1.44536e-06 $X=1500 $Y=660 $dt=0
M2 gnd3i! B Q gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.30162e-13 AS=2.28113e-13 PD=1.43036e-06 PS=1.41536e-06 $X=2340 $Y=660 $dt=0
M3 Q B gnd3i! gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.28113e-13 AS=2.30162e-13 PD=1.41536e-06 PS=1.43036e-06 $X=3230 $Y=660 $dt=0
M4 gnd3i! 7 Q gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=4.20212e-13 AS=2.28113e-13 PD=2.75536e-06 PS=1.41536e-06 $X=4070 $Y=660 $dt=0
M5 vdd3i! AN 7 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.998e-13 AS=6.768e-13 PD=2.595e-06 PS=3.78e-06 $X=620 $Y=2410 $dt=1
M6 9 7 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.115e-13 AS=6.998e-13 PD=1.71e-06 PS=2.595e-06 $X=1755 $Y=2410 $dt=1
M7 Q B 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.8775e-13 AS=2.115e-13 PD=1.96e-06 PS=1.71e-06 $X=2355 $Y=2410 $dt=1
M8 8 B Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.115e-13 AS=3.8775e-13 PD=1.71e-06 PS=1.96e-06 $X=3205 $Y=2410 $dt=1
M9 vdd3i! 7 8 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.3642e-12 AS=2.115e-13 PD=5.11e-06 PS=1.71e-06 $X=3805 $Y=2410 $dt=1
.ends NO2I1JI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX12                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX12 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=28
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=4.148e-13 AS=3.84e-13 PD=1.98e-06 PS=2.56e-06 $X=620 $Y=750 $dt=0
M1 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=4.148e-13 PD=1.34e-06 PS=1.98e-06 $X=1710 $Y=750 $dt=0
M2 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=2600 $Y=750 $dt=0
M3 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=3570 $Y=750 $dt=0
M4 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=4460 $Y=750 $dt=0
M5 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=5430 $Y=750 $dt=0
M6 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=6320 $Y=750 $dt=0
M7 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=7290 $Y=750 $dt=0
M8 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=8180 $Y=750 $dt=0
M9 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=9150 $Y=750 $dt=0
M10 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.194e-13 AS=2.16e-13 PD=1.36e-06 PS=1.34e-06 $X=10040 $Y=750 $dt=0
M11 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.84e-13 AS=2.194e-13 PD=2.56e-06 PS=1.36e-06 $X=10930 $Y=750 $dt=0
M12 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=5.79287e-13 PD=1.86506e-06 PS=3.69506e-06 $X=475 $Y=2410 $dt=1
M13 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1315 $Y=2410 $dt=1
M14 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1865 $Y=2410 $dt=1
M15 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=2705 $Y=2410 $dt=1
M16 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=3255 $Y=2410 $dt=1
M17 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=4095 $Y=2410 $dt=1
M18 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=4645 $Y=2410 $dt=1
M19 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=5485 $Y=2410 $dt=1
M20 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=6035 $Y=2410 $dt=1
M21 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=6875 $Y=2410 $dt=1
M22 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=7425 $Y=2410 $dt=1
M23 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=8265 $Y=2410 $dt=1
M24 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=8815 $Y=2410 $dt=1
M25 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=9655 $Y=2410 $dt=1
M26 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=10205 $Y=2410 $dt=1
M27 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=8.53088e-13 AS=2.54913e-13 PD=4.55506e-06 PS=1.86506e-06 $X=11045 $Y=2410 $dt=1
.ends BUJI3VX12

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INJI3VX3                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INJI3VX3 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=5 EP=4 FDC=5
M0 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=7.586e-13 PD=1.43e-06 PS=3.76e-06 $X=780 $Y=660 $dt=0
M1 gnd3i! A Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=7.586e-13 AS=2.403e-13 PD=3.76e-06 PS=1.43e-06 $X=1670 $Y=660 $dt=0
M2 Q A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=6.12287e-13 PD=1.86506e-06 PS=3.78506e-06 $X=490 $Y=2410 $dt=1
M3 vdd3i! A Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.86587e-13 AS=2.54913e-13 PD=1.88506e-06 PS=1.86506e-06 $X=1330 $Y=2410 $dt=1
M4 Q A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=5.51013e-13 AS=2.86587e-13 PD=3.69506e-06 PS=1.88506e-06 $X=1880 $Y=2410 $dt=1
.ends INJI3VX3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA4JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA4JI3VX0 vdd3i! gnd3i! D Q C B A
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 11 D gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=1.2e-13 AS=7.868e-13 PD=1.1e-06 PS=3.82e-06 $X=810 $Y=750 $dt=0
M1 10 C 11 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=1.2e-13 AS=1.2e-13 PD=1.1e-06 PS=1.1e-06 $X=1460 $Y=750 $dt=0
M2 9 B 10 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=1.2e-13 AS=1.2e-13 PD=1.1e-06 PS=1.1e-06 $X=2110 $Y=750 $dt=0
M3 Q A 9 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.84e-13 AS=1.2e-13 PD=2.56e-06 PS=1.1e-06 $X=2760 $Y=750 $dt=0
M4 Q D vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=9.882e-13 PD=1.24e-06 PS=3.92e-06 $X=540 $Y=2410 $dt=1
M5 vdd3i! C Q vdd3i! pe3i L=3e-07 W=7e-07 AD=9.882e-13 AS=1.89e-13 PD=3.92e-06 PS=1.24e-06 $X=1380 $Y=2410 $dt=1
M6 Q B vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=9.882e-13 PD=1.24e-06 PS=3.92e-06 $X=2240 $Y=2410 $dt=1
M7 vdd3i! A Q vdd3i! pe3i L=3e-07 W=7e-07 AD=9.882e-13 AS=1.89e-13 PD=3.92e-06 PS=1.24e-06 $X=3080 $Y=2410 $dt=1
.ends NA4JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OR3JI3VX1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OR3JI3VX1 vdd3i! gnd3i! A B C Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 gnd3i! A 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.482e-13 AS=2.016e-13 PD=2.04e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 8 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.116e-13 AS=2.482e-13 PD=1.78e-06 PS=2.04e-06 $X=1390 $Y=1310 $dt=0
M2 gnd3i! C 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.66689e-13 AS=2.116e-13 PD=1.17398e-06 PS=1.78e-06 $X=2160 $Y=1130 $dt=0
M3 Q 8 gnd3i! gnd3i! ne3i L=3.50112e-07 W=8.98284e-07 AD=4.174e-13 AS=3.56511e-13 PD=2.72828e-06 PS=2.51087e-06 $X=2970 $Y=660 $dt=0
M4 10 A 8 vdd3i! pe3i L=3e-07 W=1e-06 AD=1.375e-13 AS=4.8e-13 PD=1.275e-06 PS=2.96e-06 $X=670 $Y=2720 $dt=1
M5 9 B 10 vdd3i! pe3i L=3e-07 W=1e-06 AD=1.375e-13 AS=1.375e-13 PD=1.275e-06 PS=1.275e-06 $X=1245 $Y=2720 $dt=1
M6 vdd3i! C 9 vdd3i! pe3i L=3e-07 W=1e-06 AD=5.59502e-13 AS=1.375e-13 PD=2.19087e-06 PS=1.275e-06 $X=1820 $Y=2720 $dt=1
M7 Q 8 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=7.88898e-13 PD=3.78e-06 PS=3.08913e-06 $X=3000 $Y=2410 $dt=1
.ends OR3JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO3JI3VX1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO3JI3VX1 vdd3i! gnd3i! C Q B A
*.DEVICECLIMB
** N=9 EP=6 FDC=6
M0 Q C gnd3i! gnd3i! ne3i L=3.4986e-07 W=8.92071e-07 AD=2.37813e-13 AS=4.30337e-13 PD=1.42707e-06 PS=2.76707e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! B Q gnd3i! ne3i L=3.4986e-07 W=8.92071e-07 AD=2.40287e-13 AS=2.37813e-13 PD=1.44207e-06 PS=1.42707e-06 $X=1500 $Y=660 $dt=0
M2 Q A gnd3i! gnd3i! ne3i L=3.4986e-07 W=8.92071e-07 AD=4.29162e-13 AS=2.40287e-13 PD=2.74707e-06 PS=1.44207e-06 $X=2390 $Y=660 $dt=0
M3 9 C vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=1.3994e-12 PD=1.72e-06 PS=5.15e-06 $X=955 $Y=2410 $dt=1
M4 8 B 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=2.1855e-13 PD=1.72e-06 PS=1.72e-06 $X=1565 $Y=2410 $dt=1
M5 Q A 8 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=2.1855e-13 PD=3.78e-06 PS=1.72e-06 $X=2175 $Y=2410 $dt=1
.ends NO3JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: FAJI3VX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt FAJI3VX1 vdd3i! gnd3i! S CI B A CO
*.DEVICECLIMB
** N=20 EP=7 FDC=28
M0 gnd3i! 12 S gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.361e-13 AS=4.272e-13 PD=2.76e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 15 CI 12 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=7.375e-14 AS=2.832e-13 PD=8.4e-07 PS=2.14e-06 $X=2220 $Y=960 $dt=0
M2 14 B 15 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=7.375e-14 AS=7.375e-14 PD=8.4e-07 PS=8.4e-07 $X=2820 $Y=960 $dt=0
M3 gnd3i! A 14 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=2.34033e-13 AS=7.375e-14 PD=1.52158e-06 PS=8.4e-07 $X=3420 $Y=960 $dt=0
M4 13 CI gnd3i! gnd3i! ne3i L=3.5e-07 W=5.5e-07 AD=1.485e-13 AS=2.18167e-13 PD=1.09e-06 PS=1.41842e-06 $X=4350 $Y=660 $dt=0
M5 gnd3i! A 13 gnd3i! ne3i L=3.5e-07 W=5.5e-07 AD=2.5017e-13 AS=1.485e-13 PD=1.58058e-06 PS=1.09e-06 $X=5240 $Y=660 $dt=0
M6 13 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=1.296e-13 AS=2.1833e-13 PD=1.02e-06 PS=1.37942e-06 $X=6220 $Y=960 $dt=0
M7 12 10 13 gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=2.304e-13 AS=1.296e-13 PD=1.92e-06 PS=1.02e-06 $X=7110 $Y=960 $dt=0
M8 gnd3i! 10 CO gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=3.345e-13 AS=2.832e-13 PD=1.73e-06 PS=2.14e-06 $X=8700 $Y=960 $dt=0
M9 11 A gnd3i! gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=7.375e-14 AS=3.345e-13 PD=8.4e-07 PS=1.73e-06 $X=9830 $Y=960 $dt=0
M10 10 B 11 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=1.593e-13 AS=7.375e-14 PD=1.13e-06 PS=8.4e-07 $X=10430 $Y=960 $dt=0
M11 9 CI 10 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=1.593e-13 AS=1.593e-13 PD=1.13e-06 PS=1.13e-06 $X=11320 $Y=960 $dt=0
M12 gnd3i! B 9 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=4.382e-13 AS=1.593e-13 PD=1.95e-06 PS=1.13e-06 $X=12210 $Y=960 $dt=0
M13 9 A gnd3i! gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=3.068e-13 AS=4.382e-13 PD=2.22e-06 PS=1.95e-06 $X=13550 $Y=960 $dt=0
M14 vdd3i! 12 S vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.6395e-13 AS=7.1205e-13 PD=4.52213e-06 PS=3.83e-06 $X=645 $Y=2410 $dt=1
M15 vdd3i! CI 17 vdd3i! pe3i L=3e-07 W=1.03e-06 AD=4.8155e-13 AS=4.79437e-13 PD=2.35e-06 PS=3.03778e-06 $X=2125 $Y=2490 $dt=1
M16 17 B vdd3i! vdd3i! pe3i L=3e-07 W=1.03e-06 AD=3.0385e-13 AS=4.8155e-13 PD=1.62e-06 PS=2.35e-06 $X=3095 $Y=2490 $dt=1
M17 vdd3i! A 17 vdd3i! pe3i L=3e-07 W=1.03e-06 AD=4.1015e-13 AS=3.0385e-13 PD=2.01e-06 PS=1.62e-06 $X=3985 $Y=2490 $dt=1
M18 20 A vdd3i! vdd3i! pe3i L=3e-07 W=1.03e-06 AD=1.545e-13 AS=4.1015e-13 PD=1.33e-06 PS=2.01e-06 $X=4955 $Y=2490 $dt=1
M19 19 B 20 vdd3i! pe3i L=3e-07 W=1.03e-06 AD=1.545e-13 AS=1.545e-13 PD=1.33e-06 PS=1.33e-06 $X=5555 $Y=2490 $dt=1
M20 12 CI 19 vdd3i! pe3i L=3e-07 W=1.03e-06 AD=3.0385e-13 AS=1.545e-13 PD=1.62e-06 PS=1.33e-06 $X=6155 $Y=2490 $dt=1
M21 17 10 12 vdd3i! pe3i L=3e-07 W=1.03e-06 AD=6.9155e-13 AS=3.0385e-13 PD=3.77e-06 PS=1.62e-06 $X=7045 $Y=2490 $dt=1
M22 vdd3i! 10 CO vdd3i! pe3i L=3e-07 W=1.11e-06 AD=4.54624e-13 AS=5.6055e-13 PD=2.27286e-06 PS=3.23e-06 $X=8675 $Y=2410 $dt=1
M23 16 A vdd3i! vdd3i! pe3i L=3e-07 W=9.9e-07 AD=2.9205e-13 AS=4.05476e-13 PD=1.58e-06 PS=2.02714e-06 $X=9645 $Y=2530 $dt=1
M24 vdd3i! B 16 vdd3i! pe3i L=3e-07 W=9.9e-07 AD=5.763e-13 AS=2.9205e-13 PD=3.59e-06 PS=1.58e-06 $X=10535 $Y=2530 $dt=1
M25 10 CI 16 vdd3i! pe3i L=3e-07 W=1e-06 AD=2.95e-13 AS=4.65e-13 PD=1.59e-06 PS=3.01e-06 $X=12085 $Y=2520 $dt=1
M26 18 B 10 vdd3i! pe3i L=3e-07 W=1e-06 AD=1.5e-13 AS=2.95e-13 PD=1.3e-06 PS=1.59e-06 $X=12975 $Y=2520 $dt=1
M27 vdd3i! A 18 vdd3i! pe3i L=3e-07 W=1e-06 AD=8.18e-13 AS=1.5e-13 PD=4.39e-06 PS=1.3e-06 $X=13575 $Y=2520 $dt=1
.ends FAJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX4                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX4 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=11
M0 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=5.95e-07 AD=1.6065e-13 AS=5.803e-13 PD=1.135e-06 PS=3.52e-06 $X=660 $Y=955 $dt=0
M1 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=5.95e-07 AD=3.92379e-13 AS=1.6065e-13 PD=1.69084e-06 PS=1.135e-06 $X=1550 $Y=955 $dt=0
M2 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=5.86921e-13 PD=1.43e-06 PS=2.52916e-06 $X=2770 $Y=660 $dt=0
M3 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=3660 $Y=660 $dt=0
M4 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=3.494e-13 PD=2.74e-06 PS=1.86e-06 $X=4630 $Y=660 $dt=0
M5 6 A vdd3i! vdd3i! pe3i L=3e-07 W=1.1e-06 AD=2.97e-13 AS=9.042e-13 PD=1.64e-06 PS=4.66e-06 $X=710 $Y=2410 $dt=1
M6 vdd3i! A 6 vdd3i! pe3i L=3e-07 W=1.1e-06 AD=4.45401e-13 AS=2.97e-13 PD=2.09699e-06 PS=1.64e-06 $X=1550 $Y=2410 $dt=1
M7 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=5.91049e-13 PD=1.87971e-06 PS=2.78272e-06 $X=2445 $Y=2410 $dt=1
M8 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=3.3675e-13 AS=2.751e-13 PD=1.92971e-06 PS=1.87971e-06 $X=3285 $Y=2410 $dt=1
M9 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=3.3675e-13 PD=1.87971e-06 PS=1.92971e-06 $X=3935 $Y=2410 $dt=1
M10 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=6.3285e-13 AS=2.751e-13 PD=3.75971e-06 PS=1.87971e-06 $X=4775 $Y=2410 $dt=1
.ends BUJI3VX4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INJI3VX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INJI3VX1 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=5 EP=4 FDC=2
M0 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=6e-07 AD=2.88e-13 AS=6.428e-13 PD=2.16e-06 PS=3.62e-06 $X=710 $Y=950 $dt=0
M1 Q A vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=1.0562e-12 PD=3.78e-06 PS=4.76e-06 $X=760 $Y=2410 $dt=1
.ends INJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DLY2JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DLY2JI3VX1 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=12 EP=4 FDC=12
M0 gnd3i! A 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.577e-13 AS=2.016e-13 PD=1.79e-06 PS=1.8e-06 $X=620 $Y=660 $dt=0
M1 8 10 gnd3i! gnd3i! ne3i L=8e-07 W=4.2e-07 AD=2.548e-13 AS=3.577e-13 PD=1.7e-06 PS=1.79e-06 $X=1990 $Y=660 $dt=0
M2 8 10 9 gnd3i! ne3i L=8e-07 W=4.2e-07 AD=2.548e-13 AS=2.016e-13 PD=1.7e-06 PS=1.8e-06 $X=1990 $Y=1360 $dt=0
M3 gnd3i! 9 7 gnd3i! ne3i L=1e-06 W=4.2e-07 AD=3.42444e-13 AS=2.1e-13 PD=1.66718e-06 PS=1.62e-06 $X=3950 $Y=660 $dt=0
M4 6 9 7 gnd3i! ne3i L=1e-06 W=4.2e-07 AD=2.10588e-13 AS=2.1e-13 PD=1.81778e-06 PS=1.62e-06 $X=3950 $Y=1360 $dt=0
M5 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=7.25656e-13 PD=2.74e-06 PS=3.53282e-06 $X=6310 $Y=660 $dt=0
M6 vdd3i! A 10 vdd3i! pe3i L=3e-07 W=7e-07 AD=5.42937e-13 AS=3.535e-13 PD=2.69375e-06 PS=2.41e-06 $X=645 $Y=3120 $dt=1
M7 12 10 9 vdd3i! pe3i L=7.4e-07 W=4.2e-07 AD=2.8095e-13 AS=2.0035e-13 PD=1.785e-06 PS=1.77071e-06 $X=2050 $Y=2640 $dt=1
M8 12 10 vdd3i! vdd3i! pe3i L=7.4e-07 W=4.2e-07 AD=2.8095e-13 AS=3.25762e-13 PD=1.785e-06 PS=1.61625e-06 $X=2050 $Y=3400 $dt=1
M9 6 9 11 vdd3i! pe3i L=1e-06 W=4.2e-07 AD=2.856e-13 AS=2.479e-13 PD=2.2e-06 PS=1.715e-06 $X=4030 $Y=2660 $dt=1
M10 vdd3i! 9 11 vdd3i! pe3i L=1e-06 W=4.2e-07 AD=2.62018e-13 AS=2.479e-13 PD=1.40689e-06 PS=1.715e-06 $X=4030 $Y=3400 $dt=1
M11 Q 6 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.1205e-13 AS=8.79632e-13 PD=3.83e-06 PS=4.72311e-06 $X=6335 $Y=2410 $dt=1
.ends DLY2JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: SDFRRQJI3VX1                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt SDFRRQJI3VX1 vdd3i! gnd3i! SE SD RN D C Q
*.DEVICECLIMB
** N=31 EP=8 FDC=39
M0 gnd3i! SE 25 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.11575e-13 AS=2.016e-13 PD=1.6275e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 13 RN gnd3i! gnd3i! ne3i L=3.5e-07 W=5.4e-07 AD=2.079e-13 AS=2.72025e-13 PD=1.4625e-06 PS=2.0925e-06 $X=1410 $Y=660 $dt=0
M2 24 SE 13 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.617e-13 PD=6.7e-07 PS=1.1375e-06 $X=2340 $Y=960 $dt=0
M3 12 SD 24 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.163e-13 AS=5.25e-14 PD=1.45e-06 PS=6.7e-07 $X=2940 $Y=960 $dt=0
M4 23 D 12 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.163e-13 PD=6.7e-07 PS=1.45e-06 $X=3910 $Y=1000 $dt=0
M5 13 25 23 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=5.25e-14 PD=1.8e-06 PS=6.7e-07 $X=4510 $Y=1000 $dt=0
M6 gnd3i! 20 22 gnd3i! ne3i L=3.5e-07 W=7.2e-07 AD=3.01862e-13 AS=3.456e-13 PD=1.65084e-06 PS=2.4e-06 $X=6100 $Y=1090 $dt=0
M7 11 RN gnd3i! gnd3i! ne3i L=3.5e-07 W=8.85e-07 AD=2.20538e-13 AS=3.71038e-13 PD=1.77e-06 PS=2.02916e-06 $X=7070 $Y=925 $dt=0
M8 21 22 11 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.04662e-13 PD=6.7e-07 PS=8.4e-07 $X=7840 $Y=1390 $dt=0
M9 20 18 21 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=8440 $Y=1390 $dt=0
M10 12 19 20 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=1.134e-13 PD=1.8e-06 PS=9.6e-07 $X=9330 $Y=1390 $dt=0
M11 gnd3i! C 19 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.722e-13 AS=2.016e-13 PD=1.24e-06 PS=1.8e-06 $X=10920 $Y=1390 $dt=0
M12 18 19 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=1.722e-13 PD=1.8e-06 PS=1.24e-06 $X=11930 $Y=1390 $dt=0
M13 17 22 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=13520 $Y=1020 $dt=0
M14 16 18 17 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=14120 $Y=1020 $dt=0
M15 15 19 16 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=15010 $Y=1020 $dt=0
M16 10 14 15 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.47785e-13 AS=5.25e-14 PD=9.42595e-07 PS=6.7e-07 $X=15610 $Y=1020 $dt=0
M17 gnd3i! RN 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.9815e-13 AS=3.13165e-13 PD=1.56e-06 PS=1.9974e-06 $X=16540 $Y=660 $dt=0
M18 14 16 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=2.9815e-13 PD=2.74e-06 PS=1.56e-06 $X=17560 $Y=660 $dt=0
M19 Q 16 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=6.098e-13 PD=2.74e-06 PS=3.52e-06 $X=19190 $Y=660 $dt=0
M20 vdd3i! SE 25 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=5.776e-13 AS=3.456e-13 PD=2.10667e-06 PS=2.4e-06 $X=620 $Y=2800 $dt=1
M21 31 25 vdd3i! vdd3i! pe3i L=3e-07 W=9e-07 AD=1.125e-13 AS=7.22e-13 PD=1.15e-06 PS=2.63333e-06 $X=2030 $Y=2620 $dt=1
M22 28 SD 31 vdd3i! pe3i L=3e-07 W=9e-07 AD=2.43e-13 AS=1.125e-13 PD=1.44e-06 PS=1.15e-06 $X=2580 $Y=2620 $dt=1
M23 30 D 28 vdd3i! pe3i L=3e-07 W=9e-07 AD=1.125e-13 AS=2.43e-13 PD=1.15e-06 PS=1.44e-06 $X=3420 $Y=2620 $dt=1
M24 vdd3i! SE 30 vdd3i! pe3i L=3e-07 W=9e-07 AD=3.80558e-13 AS=1.125e-13 PD=1.98274e-06 PS=1.15e-06 $X=3970 $Y=2620 $dt=1
M25 22 20 vdd3i! vdd3i! pe3i L=3e-07 W=1.07e-06 AD=5.136e-13 AS=4.52442e-13 PD=3.1e-06 PS=2.35726e-06 $X=4890 $Y=2745 $dt=1
M26 vdd3i! RN 20 vdd3i! pe3i L=3e-07 W=1.02e-06 AD=9.30148e-13 AS=4.896e-13 PD=3.58417e-06 PS=3e-06 $X=6430 $Y=2800 $dt=1
M27 29 22 vdd3i! vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=3.83002e-13 PD=6.7e-07 PS=1.47583e-06 $X=7890 $Y=3060 $dt=1
M28 20 19 29 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=1.218e-13 AS=5.25e-14 PD=9.22677e-07 PS=6.7e-07 $X=8440 $Y=3060 $dt=1
M29 28 18 20 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.08e-13 AS=2.465e-13 PD=2.66e-06 PS=1.86732e-06 $X=9285 $Y=2670 $dt=1
M30 19 C vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.0675e-13 AS=6.327e-13 PD=2.37071e-06 PS=3.56e-06 $X=10970 $Y=2735 $dt=1
M31 vdd3i! 19 18 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.27981e-13 AS=4.01587e-13 PD=1.59258e-06 PS=3.03778e-06 $X=12390 $Y=2800 $dt=1
M32 27 22 vdd3i! vdd3i! pe3i L=3e-07 W=7.9e-07 AD=1.16525e-13 AS=3.59869e-13 PD=1.085e-06 PS=1.74742e-06 $X=13570 $Y=2730 $dt=1
M33 16 19 27 vdd3i! pe3i L=3e-07 W=7.9e-07 AD=2.25379e-13 AS=1.16525e-13 PD=1.73669e-06 PS=1.085e-06 $X=14165 $Y=2730 $dt=1
M34 26 18 16 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=1.19821e-13 PD=6.7e-07 PS=9.23306e-07 $X=15005 $Y=3100 $dt=1
M35 vdd3i! 14 26 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=6.29844e-13 AS=5.25e-14 PD=2.86017e-06 PS=6.7e-07 $X=15555 $Y=3100 $dt=1
M36 vdd3i! RN 16 vdd3i! pe3i L=3e-07 W=7.9e-07 AD=1.18471e-12 AS=3.19387e-13 PD=5.37983e-06 PS=2.5195e-06 $X=16775 $Y=2410 $dt=1
M37 vdd3i! 16 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=6.768e-13 PD=1.95e-06 PS=3.78e-06 $X=18400 $Y=2410 $dt=1
M38 Q 16 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=3.807e-13 PD=3.78e-06 PS=1.95e-06 $X=19240 $Y=2410 $dt=1
.ends SDFRRQJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX3                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX3 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=7
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=5.23e-13 AS=4.272e-13 PD=2.14e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.5365e-13 AS=5.23e-13 PD=1.46e-06 PS=2.14e-06 $X=1870 $Y=660 $dt=0
M2 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=7.586e-13 AS=2.5365e-13 PD=3.76e-06 PS=1.46e-06 $X=2790 $Y=660 $dt=0
M3 vdd3i! A 6 vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=6.11825e-13 AS=5.712e-13 PD=2.51971e-06 PS=3.70971e-06 $X=620 $Y=2410 $dt=1
M4 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=6.11825e-13 PD=1.87971e-06 PS=2.51971e-06 $X=1510 $Y=2410 $dt=1
M5 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=3.3675e-13 AS=2.751e-13 PD=1.92971e-06 PS=1.87971e-06 $X=2350 $Y=2410 $dt=1
M6 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=5.712e-13 AS=3.3675e-13 PD=3.70971e-06 PS=1.92971e-06 $X=3000 $Y=2410 $dt=1
.ends BUJI3VX3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INJI3VX0                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INJI3VX0 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=5 EP=4 FDC=2
M0 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=6.248e-13 PD=1.8e-06 PS=3.62e-06 $X=710 $Y=1130 $dt=0
M1 Q A vdd3i! vdd3i! pe3i L=3e-07 W=9.4e-07 AD=4.512e-13 AS=1.0092e-12 PD=2.84e-06 PS=4.76e-06 $X=760 $Y=2410 $dt=1
.ends INJI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA2JI3VX0 vdd3i! gnd3i! B Q A
*.DEVICECLIMB
** N=7 EP=5 FDC=4
M0 7 B gnd3i! gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=5.892e-13 PD=8.1e-07 PS=3.54e-06 $X=670 $Y=990 $dt=0
M1 Q A 7 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=2.688e-13 AS=7e-14 PD=2.08e-06 PS=8.1e-07 $X=1270 $Y=990 $dt=0
M2 Q B vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=1.1114e-12 PD=1.24e-06 PS=4.94e-06 $X=550 $Y=2410 $dt=1
M3 vdd3i! A Q vdd3i! pe3i L=3e-07 W=7e-07 AD=1.1114e-12 AS=1.89e-13 PD=4.94e-06 PS=1.24e-06 $X=1390 $Y=2410 $dt=1
.ends NA2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AO22JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AO22JI3VX1 vdd3i! gnd3i! B A C D Q
*.DEVICECLIMB
** N=12 EP=7 FDC=10
M0 11 B gnd3i! gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=5.768e-13 PD=8.1e-07 PS=3.52e-06 $X=660 $Y=990 $dt=0
M1 10 A 11 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=1.68e-13 AS=7e-14 PD=1.16e-06 PS=8.1e-07 $X=1260 $Y=990 $dt=0
M2 9 C 10 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=1.68e-13 PD=8.1e-07 PS=1.16e-06 $X=2210 $Y=990 $dt=0
M3 gnd3i! D 9 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=3.96017e-13 AS=7e-14 PD=1.66069e-06 PS=8.1e-07 $X=2810 $Y=990 $dt=0
M4 Q 10 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=6.29383e-13 PD=2.74e-06 PS=2.63931e-06 $X=4070 $Y=660 $dt=0
M5 vdd3i! B 12 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=2.295e-13 AS=4.868e-13 PD=1.39e-06 PS=3.75e-06 $X=460 $Y=2490 $dt=1
M6 12 A vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.868e-13 AS=2.295e-13 PD=3.75e-06 PS=1.39e-06 $X=1300 $Y=2490 $dt=1
M7 10 C 12 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=2.295e-13 AS=4.868e-13 PD=1.39e-06 PS=3.75e-06 $X=2020 $Y=2490 $dt=1
M8 12 D 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.868e-13 AS=2.295e-13 PD=3.75e-06 PS=1.39e-06 $X=2860 $Y=2490 $dt=1
M9 Q 10 vdd3i! vdd3i! pe3i L=3.01705e-07 W=1.47627e-06 AD=5.312e-13 AS=7.778e-13 PD=3.68627e-06 PS=4.46627e-06 $X=4120 $Y=2410 $dt=1
.ends AO22JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OR4JI3VX2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OR4JI3VX2 vdd3i! gnd3i! C D Q B A
*.DEVICECLIMB
** N=14 EP=7 FDC=16
M0 10 C gnd3i! gnd3i! ne3i L=3.5e-07 W=7e-07 AD=1.9155e-13 AS=3.417e-13 PD=1.255e-06 PS=2.39e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! D 10 gnd3i! ne3i L=3.5e-07 W=7e-07 AD=2.07711e-13 AS=1.9155e-13 PD=1.27673e-06 PS=1.255e-06 $X=1510 $Y=660 $dt=0
M2 12 10 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=2.64089e-13 PD=1.14e-06 PS=1.62327e-06 $X=2420 $Y=660 $dt=0
M3 Q 9 12 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=1.1125e-13 PD=1.43e-06 PS=1.14e-06 $X=3020 $Y=660 $dt=0
M4 11 9 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.2015e-13 AS=2.403e-13 PD=1.16e-06 PS=1.43e-06 $X=3910 $Y=660 $dt=0
M5 gnd3i! 10 11 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.54126e-13 AS=1.2015e-13 PD=1.60088e-06 PS=1.16e-06 $X=4530 $Y=660 $dt=0
M6 9 B gnd3i! gnd3i! ne3i L=3.5e-07 W=7e-07 AD=1.9155e-13 AS=1.99874e-13 PD=1.255e-06 PS=1.25912e-06 $X=5420 $Y=660 $dt=0
M7 gnd3i! A 9 gnd3i! ne3i L=3.5e-07 W=7e-07 AD=3.417e-13 AS=1.9155e-13 PD=2.39e-06 PS=1.255e-06 $X=6310 $Y=660 $dt=0
M8 14 C 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=6.768e-13 PD=1.66e-06 PS=3.78e-06 $X=710 $Y=2410 $dt=1
M9 vdd3i! D 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=5.47043e-13 AS=1.7625e-13 PD=2.41704e-06 PS=1.66e-06 $X=1260 $Y=2410 $dt=1
M10 Q 10 vdd3i! vdd3i! pe3i L=2.99799e-07 W=1.41828e-06 AD=3.622e-13 AS=5.50257e-13 PD=1.93828e-06 PS=2.43124e-06 $X=2210 $Y=2410 $dt=1
M11 vdd3i! 9 Q vdd3i! pe3i L=2.99799e-07 W=1.41828e-06 AD=4.987e-13 AS=3.622e-13 PD=2.36828e-06 PS=1.93828e-06 $X=3050 $Y=2410 $dt=1
M12 Q 9 vdd3i! vdd3i! pe3i L=2.99799e-07 W=1.41828e-06 AD=3.622e-13 AS=4.987e-13 PD=1.93828e-06 PS=2.36828e-06 $X=3930 $Y=2410 $dt=1
M13 vdd3i! 10 Q vdd3i! pe3i L=2.99799e-07 W=1.41828e-06 AD=5.8556e-13 AS=3.622e-13 PD=2.47136e-06 PS=1.93828e-06 $X=4770 $Y=2410 $dt=1
M14 13 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=5.8214e-13 PD=1.66e-06 PS=2.45692e-06 $X=5760 $Y=2410 $dt=1
M15 9 A 13 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=1.7625e-13 PD=3.78e-06 PS=1.66e-06 $X=6310 $Y=2410 $dt=1
.ends OR4JI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INJI3VX2                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INJI3VX2 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=5 EP=4 FDC=4
M0 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=1.296e-13 AS=4.408e-13 PD=1.02e-06 PS=3.52e-06 $X=500 $Y=1070 $dt=0
M1 gnd3i! A Q gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=4.408e-13 AS=1.296e-13 PD=3.52e-06 PS=1.02e-06 $X=1390 $Y=1070 $dt=0
M2 Q A vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=8.151e-13 PD=1.87971e-06 PS=4.50971e-06 $X=560 $Y=2410 $dt=1
M3 vdd3i! A Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=8.01e-13 AS=2.751e-13 PD=4.48971e-06 PS=1.87971e-06 $X=1400 $Y=2410 $dt=1
.ends INJI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AO21JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AO21JI3VX1 vdd3i! gnd3i! B A C Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 9 B gnd3i! gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=5.768e-13 PD=8.1e-07 PS=3.52e-06 $X=660 $Y=990 $dt=0
M1 8 A 9 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=1.708e-13 AS=7e-14 PD=1.17e-06 PS=8.1e-07 $X=1260 $Y=990 $dt=0
M2 gnd3i! C 8 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=3.94626e-13 AS=1.708e-13 PD=1.68386e-06 PS=1.17e-06 $X=2220 $Y=990 $dt=0
M3 Q 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=6.27174e-13 PD=2.74e-06 PS=2.67614e-06 $X=3510 $Y=660 $dt=0
M4 vdd3i! B 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=3.8185e-13 AS=4.08e-13 PD=2.53e-06 PS=2.66e-06 $X=620 $Y=2410 $dt=1
M5 10 A vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=2.295e-13 AS=3.8185e-13 PD=1.39e-06 PS=2.53e-06 $X=1340 $Y=2410 $dt=1
M6 8 C 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.08e-13 AS=2.295e-13 PD=2.66e-06 PS=1.39e-06 $X=2180 $Y=2410 $dt=1
M7 Q 8 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=7.0775e-13 PD=3.78e-06 PS=4.73e-06 $X=3560 $Y=2410 $dt=1
.ends AO21JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO2I1JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO2I1JI3VX1 vdd3i! gnd3i! AN Q B
*.DEVICECLIMB
** N=8 EP=5 FDC=6
M0 gnd3i! AN 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.78131e-13 AS=2.016e-13 PD=1.19267e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 Q 7 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.4285e-13 AS=3.77469e-13 PD=1.445e-06 PS=2.52733e-06 $X=1460 $Y=660 $dt=0
M2 gnd3i! B Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=6.098e-13 AS=2.4285e-13 PD=3.52e-06 PS=1.445e-06 $X=2350 $Y=660 $dt=0
M3 vdd3i! AN 7 vdd3i! pe3i L=3e-07 W=7e-07 AD=4.32009e-13 AS=3.36e-13 PD=1.71185e-06 PS=2.36e-06 $X=620 $Y=2410 $dt=1
M4 8 7 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=8.70191e-13 PD=1.66e-06 PS=3.44815e-06 $X=1740 $Y=2410 $dt=1
M5 Q B 8 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=1.7625e-13 PD=3.78e-06 PS=1.66e-06 $X=2290 $Y=2410 $dt=1
.ends NO2I1JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA3JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA3JI3VX0 vdd3i! gnd3i! C Q B A
*.DEVICECLIMB
** N=9 EP=6 FDC=6
M0 9 C gnd3i! gnd3i! ne3i L=3.5e-07 W=7e-07 AD=8.75e-14 AS=5.605e-13 PD=9.5e-07 PS=3.52e-06 $X=630 $Y=850 $dt=0
M1 8 B 9 gnd3i! ne3i L=3.5e-07 W=7e-07 AD=8.75e-14 AS=8.75e-14 PD=9.5e-07 PS=9.5e-07 $X=1230 $Y=850 $dt=0
M2 Q A 8 gnd3i! ne3i L=3.5e-07 W=7e-07 AD=3.36e-13 AS=8.75e-14 PD=2.36e-06 PS=9.5e-07 $X=1830 $Y=850 $dt=0
M3 Q C vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=5.76467e-13 PD=1.24e-06 PS=3.21333e-06 $X=470 $Y=2580 $dt=1
M4 vdd3i! B Q vdd3i! pe3i L=3e-07 W=7e-07 AD=5.76467e-13 AS=1.89e-13 PD=3.21333e-06 PS=1.24e-06 $X=1310 $Y=2580 $dt=1
M5 Q A vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=4.708e-13 AS=5.76467e-13 PD=3.92e-06 PS=3.21333e-06 $X=2040 $Y=2470 $dt=1
.ends NA3JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OR2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OR2JI3VX0 vdd3i! gnd3i! A B Q
*.DEVICECLIMB
** N=8 EP=5 FDC=6
M0 7 A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.75467e-13 PD=9.6e-07 PS=2.95333e-06 $X=530 $Y=1130 $dt=0
M1 gnd3i! B 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.75467e-13 AS=1.134e-13 PD=2.95333e-06 PS=9.6e-07 $X=1420 $Y=1130 $dt=0
M2 Q 7 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=5.75467e-13 PD=1.8e-06 PS=2.95333e-06 $X=2390 $Y=1130 $dt=0
M3 8 A 7 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=4.08e-13 PD=1.1e-06 PS=2.66e-06 $X=620 $Y=2410 $dt=1
M4 vdd3i! B 8 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=8.28174e-13 AS=1.0625e-13 PD=2.99419e-06 PS=1.1e-06 $X=1170 $Y=2410 $dt=1
M5 Q 7 vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=3.36e-13 AS=6.82026e-13 PD=2.36e-06 PS=2.46581e-06 $X=2440 $Y=2410 $dt=1
.ends OR2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AO211JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AO211JI3VX1 vdd3i! gnd3i! B A C D Q
*.DEVICECLIMB
** N=12 EP=7 FDC=10
M0 10 B gnd3i! gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=5.768e-13 PD=8.1e-07 PS=3.52e-06 $X=660 $Y=990 $dt=0
M1 9 A 10 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=1.68e-13 AS=7e-14 PD=1.16e-06 PS=8.1e-07 $X=1260 $Y=990 $dt=0
M2 gnd3i! C 9 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=3.164e-13 AS=1.68e-13 PD=1.86e-06 PS=1.16e-06 $X=2210 $Y=990 $dt=0
M3 9 D gnd3i! gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=2.464e-13 AS=3.164e-13 PD=2.08e-06 PS=1.86e-06 $X=3180 $Y=990 $dt=0
M4 Q 9 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=5.0945e-13 PD=2.74e-06 PS=3.7e-06 $X=4630 $Y=660 $dt=0
M5 vdd3i! B 12 vdd3i! pe3i L=3e-07 W=1e-06 AD=4.168e-13 AS=4.8e-13 PD=2.53e-06 PS=2.96e-06 $X=620 $Y=2410 $dt=1
M6 12 A vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.95e-13 AS=4.168e-13 PD=1.59e-06 PS=2.53e-06 $X=1410 $Y=2410 $dt=1
M7 11 C 12 vdd3i! pe3i L=3e-07 W=1e-06 AD=1.5e-13 AS=2.95e-13 PD=1.3e-06 PS=1.59e-06 $X=2300 $Y=2410 $dt=1
M8 9 D 11 vdd3i! pe3i L=3e-07 W=1e-06 AD=4.66e-13 AS=1.5e-13 PD=3.28e-06 PS=1.3e-06 $X=2900 $Y=2410 $dt=1
M9 Q 9 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=1.01495e-12 PD=3.78e-06 PS=4.82e-06 $X=4680 $Y=2410 $dt=1
.ends AO211JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: HAJI3VX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt HAJI3VX1 vdd3i! gnd3i! S B A CO
*.DEVICECLIMB
** N=12 EP=6 FDC=14
M0 gnd3i! 8 S gnd3i! ne3i L=3.49889e-07 W=8.98284e-07 AD=4.998e-13 AS=4.174e-13 PD=3.41456e-06 PS=2.72828e-06 $X=600 $Y=660 $dt=0
M1 gnd3i! A 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.52e-13 PD=1.43e-06 PS=2.74e-06 $X=2070 $Y=660 $dt=0
M2 9 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.70969e-13 AS=2.403e-13 PD=1.71986e-06 PS=1.43e-06 $X=2960 $Y=660 $dt=0
M3 8 10 9 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=3.632e-13 AS=1.79631e-13 PD=2.84284e-06 PS=1.14014e-06 $X=3850 $Y=960 $dt=0
M4 gnd3i! 10 CO gnd3i! ne3i L=3.5e-07 W=5.5e-07 AD=1.56292e-13 AS=2.4195e-13 PD=1.09236e-06 PS=2.03071e-06 $X=5380 $Y=1000 $dt=0
M5 11 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=2.52908e-13 PD=1.14e-06 PS=1.76764e-06 $X=6270 $Y=660 $dt=0
M6 10 A 11 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=1.1125e-13 PD=2.74e-06 PS=1.14e-06 $X=6870 $Y=660 $dt=0
M7 vdd3i! 8 S vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.07833e-13 AS=7.1205e-13 PD=2.97939e-06 PS=3.83e-06 $X=645 $Y=2410 $dt=1
M8 12 A vdd3i! vdd3i! pe3i L=3e-07 W=8.9e-07 AD=1.335e-13 AS=3.83667e-13 PD=1.19e-06 PS=1.88061e-06 $X=1615 $Y=2630 $dt=1
M9 8 B 12 vdd3i! pe3i L=3e-07 W=8.9e-07 AD=4.9565e-13 AS=1.335e-13 PD=2.12e-06 PS=1.19e-06 $X=2215 $Y=2630 $dt=1
M10 vdd3i! 10 8 vdd3i! pe3i L=3e-07 W=8.9e-07 AD=4.8925e-13 AS=4.9565e-13 PD=3.49e-06 PS=2.12e-06 $X=3525 $Y=2630 $dt=1
M11 vdd3i! 10 CO vdd3i! pe3i L=3e-07 W=1.11e-06 AD=4.3695e-13 AS=4.7415e-13 PD=2.09e-06 PS=3.23e-06 $X=4995 $Y=2410 $dt=1
M12 10 B vdd3i! vdd3i! pe3i L=3e-07 W=1.11e-06 AD=3.2745e-13 AS=4.3695e-13 PD=1.7e-06 PS=2.09e-06 $X=5965 $Y=2410 $dt=1
M13 vdd3i! A 10 vdd3i! pe3i L=3e-07 W=1.11e-06 AD=8.7795e-13 AS=3.2745e-13 PD=4.61e-06 PS=1.7e-06 $X=6855 $Y=2410 $dt=1
.ends HAJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OA21JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OA21JI3VX1 vdd3i! gnd3i! C A B Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 8 C 9 gnd3i! ne3i L=3.5e-07 W=5.4e-07 AD=3.313e-13 AS=2.97e-13 PD=1.95333e-06 PS=2.18e-06 $X=690 $Y=660 $dt=0
M1 8 A gnd3i! gnd3i! ne3i L=3.5e-07 W=5.4e-07 AD=3.313e-13 AS=2.592e-13 PD=1.95333e-06 PS=2.04e-06 $X=1620 $Y=1480 $dt=0
M2 gnd3i! B 8 gnd3i! ne3i L=3.5e-07 W=5.4e-07 AD=2.92808e-13 AS=3.313e-13 PD=1.47273e-06 PS=1.95333e-06 $X=2450 $Y=1010 $dt=0
M3 Q 9 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=4.82592e-13 PD=2.74e-06 PS=2.42727e-06 $X=3510 $Y=660 $dt=0
M4 9 C vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=2.295e-13 AS=1.03315e-12 PD=1.39e-06 PS=4.25e-06 $X=975 $Y=2880 $dt=1
M5 10 A 9 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=2.295e-13 PD=1.1e-06 PS=1.39e-06 $X=1815 $Y=2880 $dt=1
M6 vdd3i! B 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.77448e-13 AS=1.0625e-13 PD=1.94425e-06 PS=1.1e-06 $X=2365 $Y=2880 $dt=1
M7 Q 9 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=7.92002e-13 PD=3.78e-06 PS=3.22516e-06 $X=3560 $Y=2410 $dt=1
.ends OA21JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: EO2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt EO2JI3VX0 vdd3i! gnd3i! B A Q
*.DEVICECLIMB
** N=10 EP=5 FDC=10
M0 8 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.628e-13 PD=9.6e-07 PS=3.52e-06 $X=660 $Y=1130 $dt=0
M1 gnd3i! A 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.0445e-13 AS=1.134e-13 PD=1.34e-06 PS=9.6e-07 $X=1550 $Y=1130 $dt=0
M2 7 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.0445e-13 PD=6.7e-07 PS=1.34e-06 $X=2670 $Y=980 $dt=0
M3 Q A 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.503e-13 AS=5.25e-14 PD=1.15e-06 PS=6.7e-07 $X=3270 $Y=980 $dt=0
M4 gnd3i! 8 Q gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.0464e-12 AS=1.503e-13 PD=4.3e-06 PS=1.15e-06 $X=4200 $Y=1130 $dt=0
M5 10 B vdd3i! vdd3i! pe3i L=3e-07 W=9e-07 AD=1.35e-13 AS=7.175e-13 PD=1.2e-06 PS=4.61e-06 $X=575 $Y=2410 $dt=1
M6 8 A 10 vdd3i! pe3i L=3e-07 W=9e-07 AD=5.38188e-13 AS=1.35e-13 PD=3.13778e-06 PS=1.2e-06 $X=1175 $Y=2410 $dt=1
M7 vdd3i! B 9 vdd3i! pe3i L=3e-07 W=1.3e-06 AD=5.321e-13 AS=5.76588e-13 PD=2.43e-06 PS=3.57778e-06 $X=2795 $Y=2520 $dt=1
M8 9 A vdd3i! vdd3i! pe3i L=3e-07 W=1.3e-06 AD=3.835e-13 AS=5.321e-13 PD=1.89e-06 PS=2.43e-06 $X=3765 $Y=2410 $dt=1
M9 Q 8 9 vdd3i! pe3i L=3e-07 W=1.3e-06 AD=6.565e-13 AS=3.835e-13 PD=3.61e-06 PS=1.89e-06 $X=4655 $Y=2410 $dt=1
.ends EO2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO3JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO3JI3VX0 vdd3i! gnd3i! C Q B A
*.DEVICECLIMB
** N=9 EP=6 FDC=6
M0 Q C gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.75467e-13 PD=9.6e-07 PS=2.95333e-06 $X=615 $Y=1130 $dt=0
M1 gnd3i! B Q gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.75467e-13 AS=1.134e-13 PD=2.95333e-06 PS=9.6e-07 $X=1505 $Y=1130 $dt=0
M2 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=5.75467e-13 PD=1.8e-06 PS=2.95333e-06 $X=2390 $Y=1130 $dt=0
M3 9 C vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=1.55e-13 AS=1.3584e-12 PD=1.31e-06 PS=5.15e-06 $X=955 $Y=2410 $dt=1
M4 8 B 9 vdd3i! pe3i L=3e-07 W=1e-06 AD=1.55e-13 AS=1.55e-13 PD=1.31e-06 PS=1.31e-06 $X=1565 $Y=2410 $dt=1
M5 Q A 8 vdd3i! pe3i L=3e-07 W=1e-06 AD=4.8e-13 AS=1.55e-13 PD=2.96e-06 PS=1.31e-06 $X=2175 $Y=2410 $dt=1
.ends NO3JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AN31JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AN31JI3VX1 vdd3i! gnd3i! A B C Q D
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 10 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.335e-13 AS=6.098e-13 PD=1.19e-06 PS=3.52e-06 $X=660 $Y=660 $dt=0
M1 9 B 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.35725e-13 AS=1.335e-13 PD=1.195e-06 PS=1.19e-06 $X=1310 $Y=660 $dt=0
M2 Q C 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.0257e-13 AS=1.35725e-13 PD=1.8043e-06 PS=1.195e-06 $X=1965 $Y=660 $dt=0
M3 gnd3i! D Q gnd3i! ne3i L=3.5e-07 W=5.75e-07 AD=5.783e-13 AS=1.9548e-13 PD=3.52e-06 PS=1.1657e-06 $X=2910 $Y=975 $dt=0
M4 11 A vdd3i! vdd3i! pe3i L=3.00061e-07 W=1.44471e-06 AD=3.0525e-13 AS=5.93475e-13 PD=1.86471e-06 PS=3.72971e-06 $X=525 $Y=2425 $dt=1
M5 vdd3i! B 11 vdd3i! pe3i L=3.00061e-07 W=1.44471e-06 AD=4.42387e-13 AS=3.0525e-13 PD=2.08971e-06 PS=1.86471e-06 $X=1365 $Y=2425 $dt=1
M6 11 C vdd3i! vdd3i! pe3i L=3.00061e-07 W=1.44471e-06 AD=2.6565e-13 AS=4.42387e-13 PD=1.86471e-06 PS=2.08971e-06 $X=2310 $Y=2425 $dt=1
M7 Q D 11 vdd3i! pe3i L=3.00061e-07 W=1.44471e-06 AD=7.2375e-13 AS=2.6565e-13 PD=3.85971e-06 PS=1.86471e-06 $X=2910 $Y=2425 $dt=1
.ends AN31JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND2JI3VX0                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND2JI3VX0 vdd3i! gnd3i! A B Q
*.DEVICECLIMB
** N=8 EP=5 FDC=6
M0 7 A 8 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=2.688e-13 PD=8.1e-07 PS=2.08e-06 $X=820 $Y=990 $dt=0
M1 gnd3i! B 7 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=3.536e-13 AS=7e-14 PD=2.12571e-06 PS=8.1e-07 $X=1420 $Y=990 $dt=0
M2 Q 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=2.652e-13 PD=1.8e-06 PS=1.59429e-06 $X=2390 $Y=1130 $dt=0
M3 8 A vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=7.276e-13 PD=1.24e-06 PS=4.56e-06 $X=580 $Y=2410 $dt=1
M4 vdd3i! B 8 vdd3i! pe3i L=3e-07 W=7e-07 AD=5.276e-13 AS=1.89e-13 PD=2.48e-06 PS=1.24e-06 $X=1420 $Y=2410 $dt=1
M5 Q 8 vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=3.36e-13 AS=5.276e-13 PD=2.36e-06 PS=2.48e-06 $X=2440 $Y=2410 $dt=1
.ends AND2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO3I1JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO3I1JI3VX1 vdd3i! gnd3i! AN Q B C
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 gnd3i! AN 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.99484e-13 AS=2.016e-13 PD=1.19267e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 Q 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=4.22716e-13 PD=1.43e-06 PS=2.52733e-06 $X=1550 $Y=660 $dt=0
M2 gnd3i! B Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=2440 $Y=660 $dt=0
M3 Q C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=3.494e-13 PD=2.74e-06 PS=1.86e-06 $X=3410 $Y=660 $dt=0
M4 vdd3i! AN 8 vdd3i! pe3i L=3e-07 W=7e-07 AD=4.49443e-13 AS=3.36e-13 PD=1.73175e-06 PS=2.36e-06 $X=620 $Y=2415 $dt=1
M5 10 8 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=9.05307e-13 PD=1.72e-06 PS=3.48825e-06 $X=1770 $Y=2410 $dt=1
M6 9 B 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=2.1855e-13 PD=1.72e-06 PS=1.72e-06 $X=2380 $Y=2410 $dt=1
M7 Q C 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=2.1855e-13 PD=3.78e-06 PS=1.72e-06 $X=2990 $Y=2410 $dt=1
.ends NO3I1JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AN211JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AN211JI3VX1 vdd3i! gnd3i! B A Q C D
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 9 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=6.47e-13 PD=1.14e-06 PS=3.58e-06 $X=690 $Y=660 $dt=0
M1 Q A 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.9785e-13 AS=1.1125e-13 PD=1.71704e-06 PS=1.14e-06 $X=1290 $Y=660 $dt=0
M2 gnd3i! C Q gnd3i! ne3i L=3.5e-07 W=6.65e-07 AD=5.036e-13 AS=2.2255e-13 PD=2.145e-06 PS=1.28296e-06 $X=2250 $Y=885 $dt=0
M3 Q D gnd3i! gnd3i! ne3i L=3.5e-07 W=6.65e-07 AD=3.22525e-13 AS=5.036e-13 PD=2.3e-06 PS=2.145e-06 $X=3505 $Y=885 $dt=0
M4 vdd3i! B 11 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.5825e-13 AS=6.768e-13 PD=2.06e-06 PS=3.78e-06 $X=620 $Y=2410 $dt=1
M5 11 A vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=4.5825e-13 PD=2e-06 PS=2.06e-06 $X=1570 $Y=2410 $dt=1
M6 10 C 11 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.115e-13 AS=4.1595e-13 PD=1.71e-06 PS=2e-06 $X=2460 $Y=2410 $dt=1
M7 Q D 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=2.115e-13 PD=3.78e-06 PS=1.71e-06 $X=3060 $Y=2410 $dt=1
.ends AN211JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO22JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO22JI3VX1 vdd3i! gnd3i! B A Q C
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 8 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=4.87734e-13 PD=9.6e-07 PS=2.24324e-06 $X=720 $Y=1130 $dt=0
M1 gnd3i! A 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=4.87734e-13 AS=1.134e-13 PD=2.24324e-06 PS=9.6e-07 $X=1610 $Y=1130 $dt=0
M2 Q 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=1.03353e-12 PD=1.43e-06 PS=4.75353e-06 $X=2580 $Y=660 $dt=0
M3 gnd3i! C Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=6.098e-13 AS=2.403e-13 PD=3.52e-06 PS=1.43e-06 $X=3470 $Y=660 $dt=0
M4 10 B vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=1.0178e-12 PD=1.1e-06 PS=4.78e-06 $X=770 $Y=2410 $dt=1
M5 8 A 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.505e-13 AS=1.0625e-13 PD=2.76e-06 PS=1.1e-06 $X=1320 $Y=2410 $dt=1
M6 9 8 Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=6.768e-13 PD=1.66e-06 PS=3.78e-06 $X=2920 $Y=2410 $dt=1
M7 vdd3i! C 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=9.682e-13 AS=1.7625e-13 PD=4.66e-06 PS=1.66e-06 $X=3470 $Y=2410 $dt=1
.ends NO22JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA2JI3VX2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA2JI3VX2 vdd3i! gnd3i! B Q A
*.DEVICECLIMB
** N=8 EP=5 FDC=8
M0 8 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=7.09e-13 PD=1.14e-06 PS=3.68e-06 $X=740 $Y=660 $dt=0
M1 Q A 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=1.1125e-13 PD=1.43e-06 PS=1.14e-06 $X=1340 $Y=660 $dt=0
M2 7 A Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=2.403e-13 PD=1.14e-06 PS=1.43e-06 $X=2230 $Y=660 $dt=0
M3 gnd3i! B 7 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=7.09e-13 AS=1.1125e-13 PD=3.68e-06 PS=1.14e-06 $X=2830 $Y=660 $dt=0
M4 Q B vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.7e-13 AS=8.172e-13 PD=1.54e-06 PS=4.22e-06 $X=540 $Y=2410 $dt=1
M5 vdd3i! A Q vdd3i! pe3i L=3e-07 W=1e-06 AD=8.172e-13 AS=2.7e-13 PD=4.22e-06 PS=1.54e-06 $X=1380 $Y=2410 $dt=1
M6 Q A vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.7e-13 AS=8.172e-13 PD=1.54e-06 PS=4.22e-06 $X=2240 $Y=2410 $dt=1
M7 vdd3i! B Q vdd3i! pe3i L=3e-07 W=1e-06 AD=8.172e-13 AS=2.7e-13 PD=4.22e-06 PS=1.54e-06 $X=3080 $Y=2410 $dt=1
.ends NA2JI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO2JI3VX2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO2JI3VX2 vdd3i! gnd3i! B A Q
*.DEVICECLIMB
** N=8 EP=5 FDC=8
M0 Q B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=6.842e-13 PD=1.43e-06 PS=3.64e-06 $X=720 $Y=660 $dt=0
M1 gnd3i! A Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=1610 $Y=660 $dt=0
M2 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=2580 $Y=660 $dt=0
M3 gnd3i! B Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=6.098e-13 AS=2.403e-13 PD=3.52e-06 PS=1.43e-06 $X=3470 $Y=660 $dt=0
M4 8 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=1.6898e-12 PD=1.66e-06 PS=5.48e-06 $X=1120 $Y=2410 $dt=1
M5 Q A 8 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=1.7625e-13 PD=1.95e-06 PS=1.66e-06 $X=1670 $Y=2410 $dt=1
M6 7 A Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=3.807e-13 PD=1.66e-06 PS=1.95e-06 $X=2510 $Y=2410 $dt=1
M7 vdd3i! B 7 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.6898e-12 AS=1.7625e-13 PD=5.48e-06 PS=1.66e-06 $X=3060 $Y=2410 $dt=1
.ends NO2JI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA2I1JI3VX2                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA2I1JI3VX2 vdd3i! gnd3i! AN Q B
*.DEVICECLIMB
** N=9 EP=5 FDC=10
M0 gnd3i! AN 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.672e-13 AS=4.272e-13 PD=2.05e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 8 9 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=4.672e-13 PD=1.14e-06 PS=2.05e-06 $X=1780 $Y=660 $dt=0
M2 Q B 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.759e-13 AS=1.1125e-13 PD=1.51e-06 PS=1.14e-06 $X=2380 $Y=660 $dt=0
M3 7 B Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=2.759e-13 PD=1.14e-06 PS=1.51e-06 $X=3350 $Y=660 $dt=0
M4 gnd3i! 9 7 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=7.09e-13 AS=1.1125e-13 PD=3.68e-06 PS=1.14e-06 $X=3950 $Y=660 $dt=0
M5 vdd3i! AN 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=9.9878e-13 AS=6.768e-13 PD=4.57664e-06 PS=3.78e-06 $X=620 $Y=2410 $dt=1
M6 Q 9 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.7e-13 AS=7.08355e-13 PD=1.54e-06 PS=3.24584e-06 $X=1540 $Y=2410 $dt=1
M7 vdd3i! B Q vdd3i! pe3i L=3e-07 W=1e-06 AD=7.08355e-13 AS=2.7e-13 PD=3.24584e-06 PS=1.54e-06 $X=2380 $Y=2410 $dt=1
M8 Q B vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.7e-13 AS=7.08355e-13 PD=1.54e-06 PS=3.24584e-06 $X=3280 $Y=2410 $dt=1
M9 vdd3i! 9 Q vdd3i! pe3i L=3e-07 W=1e-06 AD=7.08355e-13 AS=2.7e-13 PD=3.24584e-06 PS=1.54e-06 $X=4120 $Y=2410 $dt=1
.ends NA2I1JI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP25JI3V                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP25JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=12
M0 gnd3i! 5 4 gnd3i! ne3i L=3.5e-07 W=8.8e-07 AD=2.376e-13 AS=4.224e-13 PD=1.42e-06 PS=2.72e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=1510 $Y=660 $dt=0
M2 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=3990 $Y=660 $dt=0
M3 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=6470 $Y=660 $dt=0
M4 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=8950 $Y=660 $dt=0
M5 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=4.312e-13 AS=2.376e-13 PD=2.74e-06 PS=1.42e-06 $X=11430 $Y=660 $dt=0
M6 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.5505e-13 AS=6.312e-13 PD=1.855e-06 PS=3.59e-06 $X=620 $Y=2505 $dt=1
M7 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.5505e-13 AS=3.5505e-13 PD=1.855e-06 PS=1.855e-06 $X=3090 $Y=2505 $dt=1
M8 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.5505e-13 AS=3.5505e-13 PD=1.855e-06 PS=1.855e-06 $X=5560 $Y=2505 $dt=1
M9 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.5505e-13 AS=3.5505e-13 PD=1.855e-06 PS=1.855e-06 $X=8030 $Y=2505 $dt=1
M10 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.84638e-13 AS=3.5505e-13 PD=1.9e-06 PS=1.855e-06 $X=10500 $Y=2505 $dt=1
M11 5 4 vdd3i! vdd3i! pe3i L=3e-07 W=1.315e-06 AD=7.56575e-13 AS=3.84638e-13 PD=3.91e-06 PS=1.9e-06 $X=13015 $Y=2505 $dt=1
.ends DECAP25JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP10JI3V                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP10JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=6
M0 gnd3i! 5 4 gnd3i! ne3i L=3.5e-07 W=8.8e-07 AD=2.376e-13 AS=4.224e-13 PD=1.42e-06 PS=2.72e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.445e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=1510 $Y=660 $dt=0
M2 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.445e-06 W=8.8e-07 AD=6.046e-13 AS=2.376e-13 PD=3.5e-06 PS=1.42e-06 $X=3495 $Y=660 $dt=0
M3 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.425e-06 W=1.315e-06 AD=3.5505e-13 AS=8.308e-13 PD=1.855e-06 PS=4.37e-06 $X=660 $Y=2505 $dt=1
M4 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.425e-06 W=1.315e-06 AD=3.71488e-13 AS=3.5505e-13 PD=1.88e-06 PS=1.855e-06 $X=2625 $Y=2505 $dt=1
M5 5 4 vdd3i! vdd3i! pe3i L=3e-07 W=1.315e-06 AD=7.56575e-13 AS=3.71488e-13 PD=3.91e-06 PS=1.88e-06 $X=4615 $Y=2505 $dt=1
.ends DECAP10JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP7JI3V                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP7JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=4
M0 gnd3i! 5 4 gnd3i! ne3i L=3.5e-07 W=8.8e-07 AD=2.376e-13 AS=4.224e-13 PD=1.42e-06 PS=2.72e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.75e-06 W=8.8e-07 AD=6.046e-13 AS=2.376e-13 PD=3.5e-06 PS=1.42e-06 $X=1510 $Y=660 $dt=0
M2 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.71e-06 W=1.315e-06 AD=3.87925e-13 AS=8.308e-13 PD=1.905e-06 PS=4.37e-06 $X=660 $Y=2505 $dt=1
M3 5 4 vdd3i! vdd3i! pe3i L=3e-07 W=1.315e-06 AD=7.237e-13 AS=3.87925e-13 PD=3.86e-06 PS=1.905e-06 $X=2960 $Y=2505 $dt=1
.ends DECAP7JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP5JI3V                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP5JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=2
M0 gnd3i! 5 4 gnd3i! ne3i L=1.48e-06 W=8.3e-07 AD=5.786e-13 AS=4.568e-13 PD=3.4e-06 PS=2.82e-06 $X=660 $Y=660 $dt=0
M1 5 4 vdd3i! vdd3i! pe3i L=1.46e-06 W=1.36e-06 AD=7.564e-13 AS=8.542e-13 PD=3.9e-06 PS=4.46e-06 $X=660 $Y=2460 $dt=1
.ends DECAP5JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP15JI3V                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP15JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=8
M0 gnd3i! 5 4 gnd3i! ne3i L=3.5e-07 W=8.8e-07 AD=2.42e-13 AS=4.224e-13 PD=1.43e-06 PS=2.72e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.71e-06 W=8.8e-07 AD=2.42e-13 AS=2.42e-13 PD=1.43e-06 PS=1.43e-06 $X=1520 $Y=660 $dt=0
M2 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.71e-06 W=8.8e-07 AD=2.376e-13 AS=2.42e-13 PD=1.42e-06 PS=1.43e-06 $X=3780 $Y=660 $dt=0
M3 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.71e-06 W=8.8e-07 AD=6.046e-13 AS=2.376e-13 PD=3.5e-06 PS=1.42e-06 $X=6030 $Y=660 $dt=0
M4 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.7e-06 W=1.315e-06 AD=3.5505e-13 AS=8.308e-13 PD=1.855e-06 PS=4.37e-06 $X=660 $Y=2505 $dt=1
M5 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.7e-06 W=1.315e-06 AD=3.5505e-13 AS=3.5505e-13 PD=1.855e-06 PS=1.855e-06 $X=2900 $Y=2505 $dt=1
M6 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.7e-06 W=1.315e-06 AD=3.78063e-13 AS=3.5505e-13 PD=1.89e-06 PS=1.855e-06 $X=5140 $Y=2505 $dt=1
M7 5 4 vdd3i! vdd3i! pe3i L=3e-07 W=1.315e-06 AD=7.56575e-13 AS=3.78063e-13 PD=3.91e-06 PS=1.89e-06 $X=7415 $Y=2505 $dt=1
.ends DECAP15JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: aska_dig                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt aska_dig 1 2 pulse_active enable DAC<5> DAC<4> DAC<3> DAC<2> DAC<1> DAC<0>
+ down_switches<21> down_switches<23> down_switches<20> down_switches<22> down_switches<19> down_switches<18> down_switches<17> down_switches<16> SPI_CS down_switches<15>
+ down_switches<13> down_switches<14> down_switches<24> porborn reset_l down_switches<27> down_switches<26> down_switches<25> down_switches<29> down_switches<30>
+ up_switches<31> up_switches<30> down_switches<28> SPI_MOSI IC_addr<1> up_switches<29> IC_addr<0> up_switches<28> up_switches<27> down_switches<31>
+ up_switches<26> up_switches<25> down_switches<12> up_switches<24> clk down_switches<2> up_switches<23> up_switches<22> down_switches<3> up_switches<21>
+ down_switches<0> up_switches<20> up_switches<19> up_switches<18> down_switches<11> up_switches<17> up_switches<16> SPI_Clk up_switches<15> up_switches<14>
+ down_switches<4> down_switches<1> down_switches<10> up_switches<13> down_switches<5> up_switches<12> down_switches<9> up_switches<11> up_switches<10> up_switches<9>
+ down_switches<8> up_switches<8> up_switches<7> up_switches<6> up_switches<5> down_switches<7> down_switches<6> up_switches<4> up_switches<3> up_switches<2>
+ up_switches<1> up_switches<0>
** N=1450 EP=82 FDC=26859
X8323 1 2 145 142 BUJI3VX2 $T=174160 87360 1 0 $X=173730 $Y=82240
X8324 1 2 612 up_switches<31> BUJI3VX2 $T=246960 24640 0 180 $X=243170 $Y=19520
X8325 1 2 1130 up_switches<30> BUJI3VX2 $T=250320 24640 0 180 $X=246530 $Y=19520
X8326 1 2 1251 up_switches<29> BUJI3VX2 $T=250880 24640 1 0 $X=250450 $Y=19520
X8327 1 2 620 568 BUJI3VX2 $T=252560 159040 0 0 $X=252130 $Y=158400
X8328 1 2 996 up_switches<28> BUJI3VX2 $T=254240 24640 1 0 $X=253810 $Y=19520
X8329 1 2 646 584 BUJI3VX2 $T=256480 203840 0 0 $X=256050 $Y=203200
X8330 1 2 177 up_switches<27> BUJI3VX2 $T=257600 24640 1 0 $X=257170 $Y=19520
X8331 1 2 613 up_switches<26> BUJI3VX2 $T=260960 24640 1 0 $X=260530 $Y=19520
X8332 1 2 617 up_switches<25> BUJI3VX2 $T=264880 24640 1 0 $X=264450 $Y=19520
X8333 1 2 180 198 BUJI3VX2 $T=266000 33600 0 0 $X=265570 $Y=32960
X8334 1 2 609 up_switches<24> BUJI3VX2 $T=268240 24640 1 0 $X=267810 $Y=19520
X8335 1 2 clk 92 BUJI3VX2 $T=273280 212800 0 180 $X=269490 $Y=207680
X8336 1 2 620 199 BUJI3VX2 $T=273840 185920 1 0 $X=273410 $Y=180800
X8337 1 2 934 up_switches<23> BUJI3VX2 $T=277760 24640 1 0 $X=277330 $Y=19520
X8338 1 2 630 up_switches<21> BUJI3VX2 $T=285040 24640 1 0 $X=284610 $Y=19520
X8339 1 2 651 up_switches<20> BUJI3VX2 $T=288960 24640 1 0 $X=288530 $Y=19520
X8340 1 2 641 up_switches<19> BUJI3VX2 $T=292320 24640 1 0 $X=291890 $Y=19520
X8341 1 2 1265 681 BUJI3VX2 $T=299040 212800 0 0 $X=298610 $Y=212160
X8342 1 2 199 219 BUJI3VX2 $T=371840 123200 0 0 $X=371410 $Y=122560
X8343 1 2 706 1040 1038 AND2JI3VX1 $T=67200 24640 1 180 $X=63410 $Y=24000
X8344 1 2 706 1217 1381 AND2JI3VX1 $T=68880 24640 0 0 $X=68450 $Y=24000
X8345 1 2 706 314 1046 AND2JI3VX1 $T=76720 33600 0 180 $X=72930 $Y=28480
X8346 1 2 706 318 1059 AND2JI3VX1 $T=84000 33600 0 180 $X=80210 $Y=28480
X8347 1 2 706 337 1063 AND2JI3VX1 $T=89040 33600 0 180 $X=85250 $Y=28480
X8348 1 2 706 852 1073 AND2JI3VX1 $T=93520 24640 0 0 $X=93090 $Y=24000
X8349 1 2 303 269 820 EN2JI3VX0 $T=70000 176960 1 180 $X=63970 $Y=176320
X8350 1 2 326 1061 1058 EN2JI3VX0 $T=84560 203840 0 180 $X=78530 $Y=198720
X8351 1 2 335 343 844 EN2JI3VX0 $T=91280 194880 1 180 $X=85250 $Y=194240
X8352 1 2 995 528 1240 EN2JI3VX0 $T=204400 194880 0 180 $X=198370 $Y=189760
X8353 1 2 1113 538 1116 EN2JI3VX0 $T=205520 212800 1 0 $X=205090 $Y=207680
X8354 1 2 642 1145 1382 EN2JI3VX0 $T=276640 221760 0 180 $X=270610 $Y=216640
X8355 1 2 965 967 964 EN2JI3VX0 $T=343280 203840 0 180 $X=337250 $Y=198720
X8356 1 2 988 1383 1299 NA2I1JI3VX1 $T=53760 203840 1 0 $X=53330 $Y=198720
X8357 1 2 1033 1035 282 NA2I1JI3VX1 $T=58800 185920 0 0 $X=58370 $Y=185280
X8358 1 2 289 282 824 NA2I1JI3VX1 $T=62160 185920 0 0 $X=61730 $Y=185280
X8359 1 2 288 102 339 NA2I1JI3VX1 $T=64960 203840 1 0 $X=64530 $Y=198720
X8360 1 2 824 273 289 NA2I1JI3VX1 $T=68880 185920 1 180 $X=65090 $Y=185280
X8361 1 2 1049 1054 1047 NA2I1JI3VX1 $T=72800 105280 1 0 $X=72370 $Y=100160
X8362 1 2 383 1047 317 NA2I1JI3VX1 $T=79520 105280 0 180 $X=75730 $Y=100160
X8363 1 2 1050 338 837 NA2I1JI3VX1 $T=77280 185920 1 0 $X=76850 $Y=180800
X8364 1 2 1045 333 326 NA2I1JI3VX1 $T=78400 194880 1 0 $X=77970 $Y=189760
X8365 1 2 326 837 1045 NA2I1JI3VX1 $T=85120 194880 0 180 $X=81330 $Y=189760
X8366 1 2 1061 342 326 NA2I1JI3VX1 $T=83440 203840 0 0 $X=83010 $Y=203200
X8367 1 2 111 1072 331 NA2I1JI3VX1 $T=94080 105280 1 180 $X=90290 $Y=104640
X8368 1 2 339 843 1071 NA2I1JI3VX1 $T=91840 203840 1 0 $X=91410 $Y=198720
X8369 1 2 854 853 127 NA2I1JI3VX1 $T=96880 185920 1 0 $X=96450 $Y=180800
X8370 1 2 357 855 1072 NA2I1JI3VX1 $T=101920 105280 1 180 $X=98130 $Y=104640
X8371 1 2 859 113 355 NA2I1JI3VX1 $T=104720 194880 0 180 $X=100930 $Y=189760
X8372 1 2 407 405 864 NA2I1JI3VX1 $T=135520 185920 1 180 $X=131730 $Y=185280
X8373 1 2 877 1088 883 NA2I1JI3VX1 $T=148960 203840 1 0 $X=148530 $Y=198720
X8374 1 2 1344 1345 473 NA2I1JI3VX1 $T=166320 203840 0 180 $X=162530 $Y=198720
X8375 1 2 538 548 1113 NA2I1JI3VX1 $T=204400 194880 0 0 $X=203970 $Y=194240
X8376 1 2 548 173 915 NA2I1JI3VX1 $T=219520 194880 1 0 $X=219090 $Y=189760
X8377 1 2 171 545 915 NA2I1JI3VX1 $T=225680 185920 1 180 $X=221890 $Y=185280
X8378 1 2 566 1121 170 NA2I1JI3VX1 $T=232400 185920 0 180 $X=228610 $Y=180800
X8379 1 2 1161 953 209 NA2I1JI3VX1 $T=313040 168000 0 0 $X=312610 $Y=167360
X8380 1 2 209 731 1161 NA2I1JI3VX1 $T=328720 168000 1 180 $X=324930 $Y=167360
X8381 1 2 956 732 209 NA2I1JI3VX1 $T=325360 194880 1 0 $X=324930 $Y=189760
X8382 1 2 967 1168 965 NA2I1JI3VX1 $T=337120 194880 0 180 $X=333330 $Y=189760
X8383 1 2 972 970 758 NA2I1JI3VX1 $T=343280 194880 1 0 $X=342850 $Y=189760
X8384 1 2 313 307 835 104 NO3I2JI3VX1 $T=78400 194880 1 180 $X=74050 $Y=194240
X8385 1 2 353 307 124 296 NO3I2JI3VX1 $T=100240 194880 0 180 $X=95890 $Y=189760
X8386 1 2 373 enable 374 1223 NO3I2JI3VX1 $T=117040 185920 0 180 $X=112690 $Y=180800
X8387 1 2 1080 307 374 425 NO3I2JI3VX1 $T=126000 194880 1 0 $X=125570 $Y=189760
X8388 1 2 1240 545 1314 1384 NO3I2JI3VX1 $T=203280 185920 1 180 $X=198930 $Y=185280
X8389 1 2 1162 966 760 959 NO3I2JI3VX1 $T=327040 176960 1 0 $X=326610 $Y=171840
X8390 1 2 reset_l 540 546 NA2JI3VX1 $T=208320 221760 1 0 $X=207890 $Y=216640
X8391 1 2 92 145 BUJI3VX1 $T=52640 24640 0 0 $X=52210 $Y=24000
X8392 1 2 699 564 BUJI3VX1 $T=66640 141120 0 0 $X=66210 $Y=140480
X8393 1 2 131 542 BUJI3VX1 $T=207200 42560 1 0 $X=206770 $Y=37440
X8394 1 2 564 921 BUJI3VX1 $T=230160 69440 0 0 $X=229730 $Y=68800
X8395 1 2 SPI_Clk 699 BUJI3VX1 $T=309120 105280 0 0 $X=308690 $Y=104640
X8396 1 2 241 1004 94 252 DFRRQJI3VX4 $T=23520 60480 1 0 $X=23090 $Y=55360
X8397 1 2 241 819 94 305 DFRRQJI3VX4 $T=59920 42560 1 0 $X=59490 $Y=37440
X8398 1 2 241 1060 94 337 DFRRQJI3VX4 $T=76720 87360 0 0 $X=76290 $Y=86720
X8399 1 2 246 1081 84 407 DFRRQJI3VX4 $T=122640 212800 1 0 $X=122210 $Y=207680
X8400 1 2 657 674 188 659 DFRRQJI3VX4 $T=302400 221760 0 180 $X=284050 $Y=216640
X8401 1 2 226 1277 184 721 DFRRQJI3VX4 $T=344400 212800 1 180 $X=326050 $Y=212160
X8402 1 2 226 1278 184 734 DFRRQJI3VX4 $T=344960 212800 0 180 $X=326610 $Y=207680
X8403 1 2 226 746 184 965 DFRRQJI3VX4 $T=355040 203840 1 180 $X=336690 $Y=203200
X8404 1 2 226 774 184 975 DFRRQJI3VX4 $T=374080 185920 0 180 $X=355730 $Y=180800
X8405 1 2 1206 1332 BUJI3VX0 $T=30240 33600 1 0 $X=29810 $Y=28480
X8406 1 2 245 1334 BUJI3VX0 $T=34160 168000 0 0 $X=33730 $Y=167360
X8407 1 2 288 1385 BUJI3VX0 $T=38640 203840 1 0 $X=38210 $Y=198720
X8408 1 2 90 254 BUJI3VX0 $T=40320 33600 0 0 $X=39890 $Y=32960
X8409 1 2 262 803 BUJI3VX0 $T=50960 168000 1 0 $X=50530 $Y=162880
X8410 1 2 260 1209 BUJI3VX0 $T=52080 203840 0 0 $X=51650 $Y=203200
X8411 1 2 318 1219 BUJI3VX0 $T=75040 96320 1 0 $X=74610 $Y=91200
X8412 1 2 1071 330 BUJI3VX0 $T=86800 203840 0 0 $X=86370 $Y=203200
X8413 1 2 852 1221 BUJI3VX0 $T=92400 96320 0 0 $X=91970 $Y=95680
X8414 1 2 426 869 BUJI3VX0 $T=140560 212800 1 0 $X=140130 $Y=207680
X8415 1 2 482 473 BUJI3VX0 $T=146160 203840 1 0 $X=145730 $Y=198720
X8416 1 2 882 883 BUJI3VX0 $T=150640 203840 0 0 $X=150210 $Y=203200
X8417 1 2 496 893 BUJI3VX0 $T=169680 221760 1 0 $X=169250 $Y=216640
X8418 1 2 638 382 BUJI3VX0 $T=185920 132160 0 180 $X=182690 $Y=127040
X8419 1 2 540 154 BUJI3VX0 $T=197120 212800 0 0 $X=196690 $Y=212160
X8420 1 2 porborn 534 BUJI3VX0 $T=205520 221760 1 0 $X=205090 $Y=216640
X8421 1 2 SPI_CS 607 BUJI3VX0 $T=218960 221760 1 0 $X=218530 $Y=216640
X8422 1 2 588 1316 BUJI3VX0 $T=243040 212800 0 0 $X=242610 $Y=212160
X8423 1 2 154 185 BUJI3VX0 $T=245840 212800 0 0 $X=245410 $Y=212160
X8424 1 2 SPI_MOSI 596 BUJI3VX0 $T=247520 221760 1 0 $X=247090 $Y=216640
X8425 1 2 686 553 BUJI3VX0 $T=250320 221760 1 0 $X=249890 $Y=216640
X8426 1 2 572 582 BUJI3VX0 $T=252000 194880 1 0 $X=251570 $Y=189760
X8427 1 2 602 604 BUJI3VX0 $T=253680 203840 0 0 $X=253250 $Y=203200
X8428 1 2 1142 1252 BUJI3VX0 $T=254800 168000 0 0 $X=254370 $Y=167360
X8429 1 2 639 930 BUJI3VX0 $T=255920 185920 1 0 $X=255490 $Y=180800
X8430 1 2 584 620 BUJI3VX0 $T=262640 176960 0 0 $X=262210 $Y=176320
X8431 1 2 584 181 BUJI3VX0 $T=263200 203840 0 0 $X=262770 $Y=203200
X8432 1 2 1382 1256 BUJI3VX0 $T=268240 221760 1 0 $X=267810 $Y=216640
X8433 1 2 621 1320 BUJI3VX0 $T=273280 185920 0 0 $X=272850 $Y=185280
X8434 1 2 190 1258 BUJI3VX0 $T=274400 176960 0 0 $X=273970 $Y=176320
X8435 1 2 638 235 BUJI3VX0 $T=277760 168000 1 0 $X=277330 $Y=162880
X8436 1 2 640 670 BUJI3VX0 $T=278320 221760 1 0 $X=277890 $Y=216640
X8437 1 2 1146 936 BUJI3VX0 $T=279440 194880 1 0 $X=279010 $Y=189760
X8438 1 2 681 646 BUJI3VX0 $T=281120 212800 0 0 $X=280690 $Y=212160
X8439 1 2 656 1148 BUJI3VX0 $T=285600 212800 1 0 $X=285170 $Y=207680
X8440 1 2 670 1265 BUJI3VX0 $T=294000 212800 1 0 $X=293570 $Y=207680
X8441 1 2 942 680 BUJI3VX0 $T=298480 194880 1 0 $X=298050 $Y=189760
X8442 1 2 1179 1285 BUJI3VX0 $T=349440 203840 1 0 $X=349010 $Y=198720
X8443 1 2 260 797 1386 288 AN21JI3VX1 $T=45360 203840 1 180 $X=41570 $Y=203200
X8444 1 2 180 798 86 257 AN21JI3VX1 $T=47040 69440 1 180 $X=43250 $Y=68800
X8445 1 2 300 813 1212 1187 AN21JI3VX1 $T=58800 194880 0 180 $X=55010 $Y=189760
X8446 1 2 131 808 274 98 AN21JI3VX1 $T=56560 42560 0 0 $X=56130 $Y=41920
X8447 1 2 102 816 313 1039 AN21JI3VX1 $T=60480 194880 0 0 $X=60050 $Y=194240
X8448 1 2 1047 108 1336 1049 AN21JI3VX1 $T=72800 105280 0 180 $X=69010 $Y=100160
X8449 1 2 343 114 850 849 AN21JI3VX1 $T=95760 185920 1 180 $X=91970 $Y=185280
X8450 1 2 1075 1072 344 357 AN21JI3VX1 $T=97440 105280 1 180 $X=93650 $Y=104640
X8451 1 2 343 1222 1387 1071 AN21JI3VX1 $T=95200 212800 0 0 $X=94770 $Y=212160
X8452 1 2 405 419 1080 130 AN21JI3VX1 $T=133280 194880 0 180 $X=129490 $Y=189760
X8453 1 2 426 412 1388 407 AN21JI3VX1 $T=136640 203840 1 180 $X=132850 $Y=203200
X8454 1 2 1305 444 1087 881 AN21JI3VX1 $T=155680 185920 0 180 $X=151890 $Y=180800
X8455 1 2 1231 425 877 420 AN21JI3VX1 $T=156800 203840 0 180 $X=153010 $Y=198720
X8456 1 2 139 425 1344 420 AN21JI3VX1 $T=162960 203840 0 180 $X=159170 $Y=198720
X8457 1 2 531 1312 1389 1314 AN21JI3VX1 $T=204400 185920 0 0 $X=203970 $Y=185280
X8458 1 2 170 1351 1390 1241 AN21JI3VX1 $T=222880 194880 1 0 $X=222450 $Y=189760
X8459 1 2 1352 159 920 558 AN21JI3VX1 $T=225680 203840 1 0 $X=225250 $Y=198720
X8460 1 2 924 925 1246 1372 AN21JI3VX1 $T=240800 185920 1 180 $X=237010 $Y=185280
X8461 1 2 734 1361 1272 721 AN21JI3VX1 $T=330960 203840 0 180 $X=327170 $Y=198720
X8462 1 2 220 724 1169 1170 AN21JI3VX1 $T=330960 185920 0 0 $X=330530 $Y=185280
X8463 1 2 1164 963 708 723 AN21JI3VX1 $T=335440 176960 1 0 $X=335010 $Y=171840
X8464 1 2 227 971 1391 969 AN21JI3VX1 $T=345520 176960 0 180 $X=341730 $Y=171840
X8465 1 2 286 88 1026 1392 EN3JI3VX1 $T=43680 96320 1 0 $X=43250 $Y=91200
X8466 1 2 1035 1187 273 1393 NA3I2JI3VX1 $T=59360 194880 1 0 $X=58930 $Y=189760
X8467 1 2 1383 1039 102 1215 NA3I2JI3VX1 $T=60480 203840 1 0 $X=60050 $Y=198720
X8468 1 2 518 514 567 167 NA3I2JI3VX1 $T=188720 194880 0 0 $X=188290 $Y=194240
X8469 1 2 1121 1241 1353 1394 NA3I2JI3VX1 $T=227360 185920 0 0 $X=226930 $Y=185280
X8470 1 2 1395 1146 642 634 NA3I2JI3VX1 $T=277760 212800 0 180 $X=273410 $Y=207680
X8471 1 2 282 1029 273 813 NA22JI3VX1 $T=54320 185920 0 0 $X=53890 $Y=185280
X8472 1 2 808 131 815 827 NA22JI3VX1 $T=61040 42560 0 0 $X=60610 $Y=41920
X8473 1 2 342 296 991 1068 NA22JI3VX1 $T=89600 203840 0 0 $X=89170 $Y=203200
X8474 1 2 440 1375 1189 419 NA22JI3VX1 $T=145600 194880 0 180 $X=141250 $Y=189760
X8475 1 2 870 876 434 460 NA22JI3VX1 $T=142240 185920 0 0 $X=141810 $Y=185280
X8476 1 2 893 420 891 499 NA22JI3VX1 $T=170800 203840 1 180 $X=166450 $Y=203200
X8477 1 2 548 159 541 558 NA22JI3VX1 $T=207760 194880 0 0 $X=207330 $Y=194240
X8478 1 2 956 708 enable 998 NA22JI3VX1 $T=313600 194880 0 0 $X=313170 $Y=194240
X8479 1 2 217 722 717 218 NA22JI3VX1 $T=333200 176960 1 180 $X=328850 $Y=176320
X8480 1 2 708 1168 enable 1274 NA22JI3VX1 $T=334880 194880 1 180 $X=330530 $Y=194240
X8481 1 2 972 708 enable 1281 NA22JI3VX1 $T=344960 194880 1 180 $X=340610 $Y=194240
X8482 1 2 1180 1330 230 749 NA22JI3VX1 $T=356160 176960 0 180 $X=351810 $Y=171840
X8483 1 2 278 801 264 804 96 AN22JI3VX1 $T=47040 51520 1 0 $X=46610 $Y=46400
X8484 1 2 1213 264 808 93 263 AN22JI3VX1 $T=56000 51520 0 180 $X=51650 $Y=46400
X8485 1 2 286 321 810 327 91 AN22JI3VX1 $T=64960 96320 1 180 $X=60610 $Y=95680
X8486 1 2 341 321 1036 327 812 AN22JI3VX1 $T=64960 105280 1 180 $X=60610 $Y=104640
X8487 1 2 276 321 821 327 100 AN22JI3VX1 $T=70000 96320 1 180 $X=65650 $Y=95680
X8488 1 2 824 1043 320 826 297 AN22JI3VX1 $T=67200 185920 1 0 $X=66770 $Y=180800
X8489 1 2 1065 112 1396 321 383 AN22JI3VX1 $T=85120 96320 1 180 $X=80770 $Y=95680
X8490 1 2 990 112 839 321 111 AN22JI3VX1 $T=90160 96320 1 180 $X=85810 $Y=95680
X8491 1 2 848 321 846 112 1303 AN22JI3VX1 $T=91280 105280 0 180 $X=86930 $Y=100160
X8492 1 2 505 353 991 124 enable AN22JI3VX1 $T=100240 194880 1 180 $X=95890 $Y=194240
X8493 1 2 876 445 878 451 452 AN22JI3VX1 $T=144480 194880 0 0 $X=144050 $Y=194240
X8494 1 2 431 151 648 180 446 AN22JI3VX1 $T=145040 24640 0 0 $X=144610 $Y=24000
X8495 1 2 1094 135 885 886 477 AN22JI3VX1 $T=160720 194880 1 180 $X=156370 $Y=194240
X8496 1 2 493 1104 480 502 1103 AN22JI3VX1 $T=176400 194880 0 180 $X=172050 $Y=189760
X8497 1 2 496 506 993 502 150 AN22JI3VX1 $T=179760 203840 1 0 $X=179330 $Y=198720
X8498 1 2 505 567 541 514 enable AN22JI3VX1 $T=184240 194880 0 0 $X=183810 $Y=194240
X8499 1 2 1246 1195 567 922 594 AN22JI3VX1 $T=236320 194880 0 180 $X=231970 $Y=189760
X8500 1 2 1260 687 776 198 940 AN22JI3VX1 $T=288400 33600 1 0 $X=287970 $Y=28480
X8501 1 2 668 687 771 198 1149 AN22JI3VX1 $T=295120 42560 0 180 $X=290770 $Y=37440
X8502 1 2 946 202 711 696 1156 AN22JI3VX1 $T=306320 168000 1 180 $X=301970 $Y=167360
X8503 1 2 1153 705 950 202 700 AN22JI3VX1 $T=304640 185920 0 0 $X=304210 $Y=185280
X8504 1 2 841 1300 DLY1JI3VX1 $T=53200 176960 1 0 $X=52770 $Y=171840
X8505 1 2 1211 275 DLY1JI3VX1 $T=53760 87360 0 0 $X=53330 $Y=86720
X8506 1 2 285 281 DLY1JI3VX1 $T=56560 69440 1 0 $X=56130 $Y=64320
X8507 1 2 291 284 DLY1JI3VX1 $T=58800 176960 1 0 $X=58370 $Y=171840
X8508 1 2 302 306 DLY1JI3VX1 $T=71120 42560 0 0 $X=70690 $Y=41920
X8509 1 2 483 834 DLY1JI3VX1 $T=73920 159040 0 0 $X=73490 $Y=158400
X8510 1 2 309 319 DLY1JI3VX1 $T=76720 51520 0 0 $X=76290 $Y=50880
X8511 1 2 1064 325 DLY1JI3VX1 $T=79520 159040 0 0 $X=79090 $Y=158400
X8512 1 2 323 328 DLY1JI3VX1 $T=82880 33600 0 0 $X=82450 $Y=32960
X8513 1 2 840 332 DLY1JI3VX1 $T=84000 176960 0 0 $X=83570 $Y=176320
X8514 1 2 384 366 DLY1JI3VX1 $T=88480 33600 0 0 $X=88050 $Y=32960
X8515 1 2 354 1367 DLY1JI3VX1 $T=89600 176960 0 0 $X=89170 $Y=176320
X8516 1 2 388 1069 DLY1JI3VX1 $T=99680 42560 1 180 $X=93650 $Y=41920
X8517 1 2 1074 1338 DLY1JI3VX1 $T=96880 24640 0 0 $X=96450 $Y=24000
X8518 1 2 362 361 DLY1JI3VX1 $T=105280 42560 1 180 $X=99250 $Y=41920
X8519 1 2 390 363 DLY1JI3VX1 $T=105280 87360 0 180 $X=99250 $Y=82240
X8520 1 2 428 857 DLY1JI3VX1 $T=105280 105280 0 180 $X=99250 $Y=100160
X8521 1 2 381 117 DLY1JI3VX1 $T=105280 150080 0 180 $X=99250 $Y=144960
X8522 1 2 385 120 DLY1JI3VX1 $T=113120 78400 1 0 $X=112690 $Y=73280
X8523 1 2 389 370 DLY1JI3VX1 $T=113120 78400 0 0 $X=112690 $Y=77760
X8524 1 2 423 371 DLY1JI3VX1 $T=113120 96320 0 0 $X=112690 $Y=95680
X8525 1 2 378 125 DLY1JI3VX1 $T=113120 150080 0 0 $X=112690 $Y=149440
X8526 1 2 387 375 DLY1JI3VX1 $T=116480 24640 0 0 $X=116050 $Y=24000
X8527 1 2 497 377 DLY1JI3VX1 $T=117600 123200 1 0 $X=117170 $Y=118080
X8528 1 2 861 862 DLY1JI3VX1 $T=118720 96320 0 0 $X=118290 $Y=95680
X8529 1 2 519 394 DLY1JI3VX1 $T=123200 123200 1 0 $X=122770 $Y=118080
X8530 1 2 128 395 DLY1JI3VX1 $T=123200 176960 0 0 $X=122770 $Y=176320
X8531 1 2 406 415 DLY1JI3VX1 $T=133840 33600 0 0 $X=133410 $Y=32960
X8532 1 2 438 416 DLY1JI3VX1 $T=133840 69440 0 0 $X=133410 $Y=68800
X8533 1 2 494 422 DLY1JI3VX1 $T=137760 114240 0 0 $X=137330 $Y=113600
X8534 1 2 526 424 DLY1JI3VX1 $T=138320 132160 0 0 $X=137890 $Y=131520
X8535 1 2 500 439 DLY1JI3VX1 $T=142800 141120 1 0 $X=142370 $Y=136000
X8536 1 2 524 441 DLY1JI3VX1 $T=143360 114240 1 0 $X=142930 $Y=109120
X8537 1 2 429 443 DLY1JI3VX1 $T=143920 51520 1 0 $X=143490 $Y=46400
X8538 1 2 1342 449 DLY1JI3VX1 $T=145040 176960 0 0 $X=144610 $Y=176320
X8539 1 2 455 880 DLY1JI3VX1 $T=145600 168000 1 0 $X=145170 $Y=162880
X8540 1 2 1230 456 DLY1JI3VX1 $T=150640 51520 1 0 $X=150210 $Y=46400
X8541 1 2 484 1190 DLY1JI3VX1 $T=150640 176960 0 0 $X=150210 $Y=176320
X8542 1 2 433 133 DLY1JI3VX1 $T=151200 168000 1 0 $X=150770 $Y=162880
X8543 1 2 1106 464 DLY1JI3VX1 $T=154000 123200 0 0 $X=153570 $Y=122560
X8544 1 2 498 465 DLY1JI3VX1 $T=154000 141120 1 0 $X=153570 $Y=136000
X8545 1 2 134 468 DLY1JI3VX1 $T=155120 150080 1 0 $X=154690 $Y=144960
X8546 1 2 459 1098 DLY1JI3VX1 $T=156240 51520 1 0 $X=155810 $Y=46400
X8547 1 2 895 1100 DLY1JI3VX1 $T=159040 168000 0 0 $X=158610 $Y=167360
X8548 1 2 469 478 DLY1JI3VX1 $T=160720 42560 1 0 $X=160290 $Y=37440
X8549 1 2 1234 892 DLY1JI3VX1 $T=164080 159040 1 0 $X=163650 $Y=153920
X8550 1 2 549 1306 DLY1JI3VX1 $T=164080 221760 1 0 $X=163650 $Y=216640
X8551 1 2 1346 894 DLY1JI3VX1 $T=166880 42560 1 0 $X=166450 $Y=37440
X8552 1 2 140 486 DLY1JI3VX1 $T=168000 78400 1 0 $X=167570 $Y=73280
X8553 1 2 479 487 DLY1JI3VX1 $T=168560 87360 1 0 $X=168130 $Y=82240
X8554 1 2 491 144 DLY1JI3VX1 $T=172480 42560 1 0 $X=172050 $Y=37440
X8555 1 2 523 158 DLY1JI3VX1 $T=183120 24640 1 180 $X=177090 $Y=24000
X8556 1 2 1237 504 DLY1JI3VX1 $T=178640 60480 1 0 $X=178210 $Y=55360
X8557 1 2 901 513 DLY1JI3VX1 $T=182560 150080 1 0 $X=182130 $Y=144960
X8558 1 2 1109 516 DLY1JI3VX1 $T=184240 194880 1 0 $X=183810 $Y=189760
X8559 1 2 1307 521 DLY1JI3VX1 $T=189280 33600 1 0 $X=188850 $Y=28480
X8560 1 2 520 522 DLY1JI3VX1 $T=189280 60480 1 0 $X=188850 $Y=55360
X8561 1 2 1308 1110 DLY1JI3VX1 $T=196000 78400 0 180 $X=189970 $Y=73280
X8562 1 2 994 905 DLY1JI3VX1 $T=194880 33600 1 0 $X=194450 $Y=28480
X8563 1 2 525 907 DLY1JI3VX1 $T=197680 141120 0 0 $X=197250 $Y=140480
X8564 1 2 155 530 DLY1JI3VX1 $T=199360 221760 1 0 $X=198930 $Y=216640
X8565 1 2 562 166 DLY1JI3VX1 $T=205520 60480 1 180 $X=199490 $Y=59840
X8566 1 2 911 156 DLY1JI3VX1 $T=203280 141120 0 0 $X=202850 $Y=140480
X8567 1 2 543 1311 DLY1JI3VX1 $T=211120 60480 1 180 $X=205090 $Y=59840
X8568 1 2 539 1363 DLY1JI3VX1 $T=211120 87360 0 180 $X=205090 $Y=82240
X8569 1 2 544 1194 DLY1JI3VX1 $T=211120 185920 0 180 $X=205090 $Y=180800
X8570 1 2 165 162 DLY1JI3VX1 $T=218960 176960 0 0 $X=218530 $Y=176320
X8571 1 2 563 164 DLY1JI3VX1 $T=225120 87360 0 180 $X=219090 $Y=82240
X8572 1 2 1244 555 DLY1JI3VX1 $T=230720 87360 0 180 $X=224690 $Y=82240
X8573 1 2 1245 163 DLY1JI3VX1 $T=235200 33600 0 180 $X=229170 $Y=28480
X8574 1 2 1124 569 DLY1JI3VX1 $T=230720 87360 1 0 $X=230290 $Y=82240
X8575 1 2 599 179 DLY1JI3VX1 $T=238000 87360 1 0 $X=237570 $Y=82240
X8576 1 2 186 590 DLY1JI3VX1 $T=240800 24640 0 0 $X=240370 $Y=24000
X8577 1 2 182 638 DLY1JI3VX1 $T=244160 168000 0 0 $X=243730 $Y=167360
X8578 1 2 587 595 DLY1JI3VX1 $T=244160 176960 1 0 $X=243730 $Y=171840
X8579 1 2 607 182 DLY1JI3VX1 $T=244720 159040 0 0 $X=244290 $Y=158400
X8580 1 2 593 600 DLY1JI3VX1 $T=248080 60480 0 0 $X=247650 $Y=59840
X8581 1 2 1250 605 DLY1JI3VX1 $T=250320 33600 1 0 $X=249890 $Y=28480
X8582 1 2 1196 187 DLY1JI3VX1 $T=251440 176960 1 0 $X=251010 $Y=171840
X8583 1 2 601 189 DLY1JI3VX1 $T=253680 60480 0 0 $X=253250 $Y=59840
X8584 1 2 1253 997 DLY1JI3VX1 $T=257040 176960 0 0 $X=256610 $Y=176320
X8585 1 2 1356 618 DLY1JI3VX1 $T=259840 42560 0 0 $X=259410 $Y=41920
X8586 1 2 649 635 DLY1JI3VX1 $T=262080 60480 0 0 $X=261650 $Y=59840
X8587 1 2 1254 191 DLY1JI3VX1 $T=265440 42560 0 0 $X=265010 $Y=41920
X8588 1 2 933 631 DLY1JI3VX1 $T=267680 176960 0 0 $X=267250 $Y=176320
X8589 1 2 629 935 DLY1JI3VX1 $T=271600 42560 0 0 $X=271170 $Y=41920
X8590 1 2 937 645 DLY1JI3VX1 $T=277200 42560 0 0 $X=276770 $Y=41920
X8591 1 2 939 652 DLY1JI3VX1 $T=282800 60480 0 0 $X=282370 $Y=59840
X8592 1 2 1259 941 DLY1JI3VX1 $T=283360 176960 0 0 $X=282930 $Y=176320
X8593 1 2 653 665 DLY1JI3VX1 $T=288400 60480 0 0 $X=287970 $Y=59840
X8594 1 2 655 667 DLY1JI3VX1 $T=288960 176960 0 0 $X=288530 $Y=176320
X8595 1 2 679 678 DLY1JI3VX1 $T=294560 60480 0 0 $X=294130 $Y=59840
X8596 1 2 1323 684 DLY1JI3VX1 $T=300160 42560 0 0 $X=299730 $Y=41920
X8597 1 2 1266 201 DLY1JI3VX1 $T=300160 60480 1 0 $X=299730 $Y=55360
X8598 1 2 185 686 DLY1JI3VX1 $T=302400 221760 1 0 $X=301970 $Y=216640
X8599 1 2 948 695 DLY1JI3VX1 $T=304080 87360 0 0 $X=303650 $Y=86720
X8600 1 2 693 1199 DLY1JI3VX1 $T=311360 60480 0 180 $X=305330 $Y=55360
X8601 1 2 685 702 DLY1JI3VX1 $T=306320 168000 0 0 $X=305890 $Y=167360
X8602 1 2 1270 707 DLY1JI3VX1 $T=309680 87360 1 0 $X=309250 $Y=82240
X8603 1 2 710 1359 DLY1JI3VX1 $T=316960 60480 0 180 $X=310930 $Y=55360
X8604 1 2 207 952 DLY1JI3VX1 $T=316960 150080 0 180 $X=310930 $Y=144960
X8605 1 2 208 1200 DLY1JI3VX1 $T=316960 150080 1 180 $X=310930 $Y=149440
X8606 1 2 726 211 DLY1JI3VX1 $T=324800 78400 0 0 $X=324370 $Y=77760
X8607 1 2 728 216 DLY1JI3VX1 $T=324800 105280 0 0 $X=324370 $Y=104640
X8608 1 2 1167 729 DLY1JI3VX1 $T=330400 51520 1 0 $X=329970 $Y=46400
X8609 1 2 1275 1174 DLY1JI3VX1 $T=334880 60480 1 0 $X=334450 $Y=55360
X8610 1 2 1380 737 DLY1JI3VX1 $T=334880 168000 1 0 $X=334450 $Y=162880
X8611 1 2 765 1201 DLY1JI3VX1 $T=340480 168000 1 0 $X=340050 $Y=162880
X8612 1 2 1327 1328 DLY1JI3VX1 $T=341040 60480 1 0 $X=340610 $Y=55360
X8613 1 2 1282 747 DLY1JI3VX1 $T=346640 60480 1 0 $X=346210 $Y=55360
X8614 1 2 1329 980 DLY1JI3VX1 $T=350000 150080 0 0 $X=349570 $Y=149440
X8615 1 2 1287 753 DLY1JI3VX1 $T=351680 42560 0 0 $X=351250 $Y=41920
X8616 1 2 762 754 DLY1JI3VX1 $T=351680 51520 1 0 $X=351250 $Y=46400
X8617 1 2 1288 756 DLY1JI3VX1 $T=352240 60480 1 0 $X=351810 $Y=55360
X8618 1 2 763 764 DLY1JI3VX1 $T=355600 150080 0 0 $X=355170 $Y=149440
X8619 1 2 984 769 DLY1JI3VX1 $T=358400 176960 0 0 $X=357970 $Y=176320
X8620 1 2 772 234 DLY1JI3VX1 $T=367360 60480 0 0 $X=366930 $Y=59840
X8621 1 2 1331 777 DLY1JI3VX1 $T=367920 51520 0 0 $X=367490 $Y=50880
X8622 1 2 985 778 DLY1JI3VX1 $T=373520 51520 0 0 $X=373090 $Y=50880
X8623 1 2 986 779 DLY1JI3VX1 $T=373520 60480 0 0 $X=373090 $Y=59840
X8624 1 2 1184 780 DLY1JI3VX1 $T=373520 176960 1 0 $X=373090 $Y=171840
X8625 1 2 236 781 DLY1JI3VX1 $T=374080 33600 1 0 $X=373650 $Y=28480
X8626 1 2 1293 787 DLY1JI3VX1 $T=379120 42560 1 0 $X=378690 $Y=37440
X8627 1 2 1295 788 DLY1JI3VX1 $T=379120 42560 0 0 $X=378690 $Y=41920
X8628 1 2 1294 789 DLY1JI3VX1 $T=379120 168000 1 0 $X=378690 $Y=162880
X8629 1 2 1397 461 1224 down_switches<21> ON21JI3VX4 $T=114800 24640 1 0 $X=114370 $Y=19520
X8630 1 2 1079 461 1227 down_switches<23> ON21JI3VX4 $T=124320 24640 1 0 $X=123890 $Y=19520
X8631 1 2 868 461 867 down_switches<20> ON21JI3VX4 $T=132720 24640 1 0 $X=132290 $Y=19520
X8632 1 2 879 461 1229 down_switches<22> ON21JI3VX4 $T=150080 24640 0 180 $X=141250 $Y=19520
X8633 1 2 875 461 992 down_switches<19> ON21JI3VX4 $T=146160 33600 1 0 $X=145730 $Y=28480
X8634 1 2 1092 461 1232 down_switches<18> ON21JI3VX4 $T=159040 24640 0 180 $X=150210 $Y=19520
X8635 1 2 1101 461 1235 down_switches<17> ON21JI3VX4 $T=168000 24640 0 180 $X=159170 $Y=19520
X8636 1 2 897 461 485 down_switches<16> ON21JI3VX4 $T=176400 24640 0 180 $X=167570 $Y=19520
X8637 1 2 1398 461 1105 down_switches<15> ON21JI3VX4 $T=182000 33600 0 180 $X=173170 $Y=28480
X8638 1 2 1399 461 1107 down_switches<14> ON21JI3VX4 $T=185360 24640 0 180 $X=176530 $Y=19520
X8639 1 2 1400 461 1369 down_switches<24> ON21JI3VX4 $T=194880 33600 1 180 $X=186050 $Y=32960
X8640 1 2 1401 461 1112 down_switches<13> ON21JI3VX4 $T=197680 24640 0 180 $X=188850 $Y=19520
X8641 1 2 914 461 1313 down_switches<26> ON21JI3VX4 $T=204400 24640 1 0 $X=203970 $Y=19520
X8642 1 2 1310 461 1115 down_switches<25> ON21JI3VX4 $T=204960 33600 1 0 $X=204530 $Y=28480
X8643 1 2 1118 461 1117 down_switches<27> ON21JI3VX4 $T=225120 33600 1 180 $X=216290 $Y=32960
X8644 1 2 1123 461 1242 down_switches<29> ON21JI3VX4 $T=228480 24640 0 180 $X=219650 $Y=19520
X8645 1 2 1402 461 1249 down_switches<30> ON21JI3VX4 $T=246960 33600 0 180 $X=238130 $Y=28480
X8646 1 2 929 461 1131 down_switches<28> ON21JI3VX4 $T=253120 33600 1 180 $X=244290 $Y=32960
X8647 1 2 1319 461 1255 down_switches<31> ON21JI3VX4 $T=270480 33600 0 180 $X=261650 $Y=28480
X8648 1 2 1257 461 1139 down_switches<12> ON21JI3VX4 $T=273840 24640 1 180 $X=265010 $Y=24000
X8649 1 2 1403 461 1321 down_switches<2> ON21JI3VX4 $T=283920 33600 0 180 $X=275090 $Y=28480
X8650 1 2 1262 461 1261 down_switches<3> ON21JI3VX4 $T=291200 33600 1 180 $X=282370 $Y=32960
X8651 1 2 944 461 1264 down_switches<0> ON21JI3VX4 $T=301840 33600 0 180 $X=293010 $Y=28480
X8652 1 2 951 461 1267 down_switches<11> ON21JI3VX4 $T=309120 24640 1 180 $X=300290 $Y=24000
X8653 1 2 1404 461 1378 down_switches<1> ON21JI3VX4 $T=310800 42560 1 0 $X=310370 $Y=37440
X8654 1 2 957 461 212 down_switches<10> ON21JI3VX4 $T=310800 42560 0 0 $X=310370 $Y=41920
X8655 1 2 1405 461 999 down_switches<4> ON21JI3VX4 $T=331520 33600 0 180 $X=322690 $Y=28480
X8656 1 2 1406 461 1379 down_switches<5> ON21JI3VX4 $T=337120 24640 0 180 $X=328290 $Y=19520
X8657 1 2 1173 461 1326 down_switches<9> ON21JI3VX4 $T=341040 33600 1 180 $X=332210 $Y=32960
X8658 1 2 979 461 1284 down_switches<8> ON21JI3VX4 $T=351680 33600 1 180 $X=342850 $Y=32960
X8659 1 2 1183 461 766 down_switches<6> ON21JI3VX4 $T=366240 24640 0 180 $X=357410 $Y=19520
X8660 1 2 1407 461 1291 down_switches<7> ON21JI3VX4 $T=367920 33600 0 180 $X=359090 $Y=28480
X8661 1 2 129 489 INJI3VX6 $T=176960 168000 1 0 $X=176530 $Y=162880
X8662 1 2 252 1408 247 1009 NA3I1JI3VX1 $T=29680 60480 0 0 $X=29250 $Y=59840
X8663 1 2 93 1409 305 254 NA3I1JI3VX1 $T=56000 33600 1 180 $X=51650 $Y=32960
X8664 1 2 131 1362 815 305 NA3I1JI3VX1 $T=70000 33600 1 180 $X=65650 $Y=32960
X8665 1 2 851 842 844 843 NA3I1JI3VX1 $T=90160 194880 0 180 $X=85810 $Y=189760
X8666 1 2 173 1122 557 159 NA3I1JI3VX1 $T=227360 194880 0 0 $X=226930 $Y=194240
X8667 1 2 1122 1410 570 582 NA3I1JI3VX1 $T=236320 203840 1 0 $X=235890 $Y=198720
X8668 1 2 669 1395 663 666 NA3I1JI3VX1 $T=283360 212800 0 180 $X=279010 $Y=207680
X8669 1 2 706 pulse_active BUJI3VX8 $T=63840 24640 1 180 $X=55010 $Y=24000
X8670 1 2 1038 DAC<5> BUJI3VX8 $T=61600 24640 1 0 $X=61170 $Y=19520
X8671 1 2 1046 DAC<4> BUJI3VX8 $T=70560 24640 1 0 $X=70130 $Y=19520
X8672 1 2 1381 DAC<3> BUJI3VX8 $T=73360 24640 0 0 $X=72930 $Y=24000
X8673 1 2 1059 DAC<2> BUJI3VX8 $T=79520 24640 1 0 $X=79090 $Y=19520
X8674 1 2 1063 DAC<1> BUJI3VX8 $T=83440 24640 0 0 $X=83010 $Y=24000
X8675 1 2 1073 DAC<0> BUJI3VX8 $T=97440 24640 0 180 $X=88610 $Y=19520
X8676 1 2 142 84 BUJI3VX8 $T=173040 168000 1 180 $X=164210 $Y=167360
X8677 1 2 142 94 BUJI3VX8 $T=182560 78400 0 180 $X=173730 $Y=73280
X8678 1 2 142 184 BUJI3VX8 $T=190400 168000 0 180 $X=181570 $Y=162880
X8679 1 2 142 178 BUJI3VX8 $T=193760 87360 1 0 $X=193330 $Y=82240
X8680 1 2 241 793 84 243 DFRRQJI3VX1 $T=24080 123200 0 0 $X=23650 $Y=122560
X8681 1 2 241 237 84 240 DFRRQJI3VX1 $T=24080 141120 1 0 $X=23650 $Y=136000
X8682 1 2 241 238 84 85 DFRRQJI3VX1 $T=24080 141120 0 0 $X=23650 $Y=140480
X8683 1 2 241 1296 94 265 DFRRQJI3VX1 $T=24640 96320 0 0 $X=24210 $Y=95680
X8684 1 2 241 248 84 258 DFRRQJI3VX1 $T=24640 159040 1 0 $X=24210 $Y=153920
X8685 1 2 241 239 84 245 DFRRQJI3VX1 $T=24640 176960 1 0 $X=24210 $Y=171840
X8686 1 2 241 1332 94 93 DFRRQJI3VX1 $T=25200 33600 0 0 $X=24770 $Y=32960
X8687 1 2 241 251 94 90 DFRRQJI3VX1 $T=25200 42560 1 0 $X=24770 $Y=37440
X8688 1 2 241 1364 94 1009 DFRRQJI3VX1 $T=25200 51520 0 0 $X=24770 $Y=50880
X8689 1 2 241 1006 94 247 DFRRQJI3VX1 $T=25200 78400 1 0 $X=24770 $Y=73280
X8690 1 2 246 249 84 279 DFRRQJI3VX1 $T=25200 185920 1 0 $X=24770 $Y=180800
X8691 1 2 246 250 84 289 DFRRQJI3VX1 $T=25200 185920 0 0 $X=24770 $Y=185280
X8692 1 2 241 1204 94 1014 DFRRQJI3VX1 $T=25760 87360 1 0 $X=25330 $Y=82240
X8693 1 2 241 242 94 88 DFRRQJI3VX1 $T=25760 96320 1 0 $X=25330 $Y=91200
X8694 1 2 246 792 84 89 DFRRQJI3VX1 $T=26320 194880 0 0 $X=25890 $Y=194240
X8695 1 2 246 1007 84 288 DFRRQJI3VX1 $T=27440 212800 1 0 $X=27010 $Y=207680
X8696 1 2 241 1018 84 91 DFRRQJI3VX1 $T=39200 132160 1 0 $X=38770 $Y=127040
X8697 1 2 241 1019 84 100 DFRRQJI3VX1 $T=39760 132160 0 0 $X=39330 $Y=131520
X8698 1 2 241 799 84 259 DFRRQJI3VX1 $T=39760 141120 1 0 $X=39330 $Y=136000
X8699 1 2 246 806 84 262 DFRRQJI3VX1 $T=54880 168000 1 180 $X=39330 $Y=167360
X8700 1 2 241 275 94 257 DFRRQJI3VX1 $T=59360 87360 0 180 $X=43810 $Y=82240
X8701 1 2 246 1335 84 260 DFRRQJI3VX1 $T=44240 212800 1 0 $X=43810 $Y=207680
X8702 1 2 246 268 84 1037 DFRRQJI3VX1 $T=45360 212800 0 0 $X=44930 $Y=212160
X8703 1 2 241 1030 94 1040 DFRRQJI3VX1 $T=48160 78400 0 0 $X=47730 $Y=77760
X8704 1 2 241 281 94 283 DFRRQJI3VX1 $T=48720 69440 0 0 $X=48290 $Y=68800
X8705 1 2 241 99 94 1217 DFRRQJI3VX1 $T=48720 78400 1 0 $X=48290 $Y=73280
X8706 1 2 241 307 84 1211 DFRRQJI3VX1 $T=68320 159040 1 180 $X=52770 $Y=158400
X8707 1 2 241 817 84 298 DFRRQJI3VX1 $T=53760 159040 1 0 $X=53330 $Y=153920
X8708 1 2 241 284 84 824 DFRRQJI3VX1 $T=53760 168000 1 0 $X=53330 $Y=162880
X8709 1 2 241 1300 84 297 DFRRQJI3VX1 $T=54880 168000 0 0 $X=54450 $Y=167360
X8710 1 2 241 1216 84 812 DFRRQJI3VX1 $T=70560 132160 0 180 $X=55010 $Y=127040
X8711 1 2 241 304 84 825 DFRRQJI3VX1 $T=55440 141120 1 0 $X=55010 $Y=136000
X8712 1 2 241 299 84 317 DFRRQJI3VX1 $T=56560 114240 1 0 $X=56130 $Y=109120
X8713 1 2 241 287 84 823 DFRRQJI3VX1 $T=56560 123200 0 0 $X=56130 $Y=122560
X8714 1 2 241 827 94 131 DFRRQJI3VX1 $T=76160 51520 0 180 $X=60610 $Y=46400
X8715 1 2 241 319 94 278 DFRRQJI3VX1 $T=76720 51520 1 180 $X=61170 $Y=50880
X8716 1 2 241 306 94 96 DFRRQJI3VX1 $T=76720 60480 0 180 $X=61170 $Y=55360
X8717 1 2 246 1041 84 308 DFRRQJI3VX1 $T=61600 212800 0 0 $X=61170 $Y=212160
X8718 1 2 246 1048 84 293 DFRRQJI3VX1 $T=76720 221760 0 180 $X=61170 $Y=216640
X8719 1 2 241 312 94 309 DFRRQJI3VX1 $T=77280 60480 1 180 $X=61730 $Y=59840
X8720 1 2 241 348 94 302 DFRRQJI3VX1 $T=77840 69440 0 180 $X=62290 $Y=64320
X8721 1 2 241 1042 94 314 DFRRQJI3VX1 $T=63840 78400 0 0 $X=63410 $Y=77760
X8722 1 2 241 1044 94 318 DFRRQJI3VX1 $T=63840 87360 1 0 $X=63410 $Y=82240
X8723 1 2 241 349 94 285 DFRRQJI3VX1 $T=79520 69440 1 180 $X=63970 $Y=68800
X8724 1 2 241 316 84 324 DFRRQJI3VX1 $T=69440 150080 0 0 $X=69010 $Y=149440
X8725 1 2 241 109 84 291 DFRRQJI3VX1 $T=84560 159040 0 180 $X=69010 $Y=153920
X8726 1 2 241 834 84 295 DFRRQJI3VX1 $T=84560 168000 0 180 $X=69010 $Y=162880
X8727 1 2 241 332 84 339 DFRRQJI3VX1 $T=84560 176960 0 180 $X=69010 $Y=171840
X8728 1 2 241 325 84 1045 DFRRQJI3VX1 $T=85120 168000 1 180 $X=69570 $Y=167360
X8729 1 2 241 328 94 376 DFRRQJI3VX1 $T=77840 42560 1 0 $X=77410 $Y=37440
X8730 1 2 241 350 94 362 DFRRQJI3VX1 $T=77840 42560 0 0 $X=77410 $Y=41920
X8731 1 2 241 107 94 323 DFRRQJI3VX1 $T=92960 51520 0 180 $X=77410 $Y=46400
X8732 1 2 246 329 84 326 DFRRQJI3VX1 $T=93520 212800 1 180 $X=77970 $Y=212160
X8733 1 2 246 1062 84 343 DFRRQJI3VX1 $T=78400 221760 1 0 $X=77970 $Y=216640
X8734 1 2 241 1066 94 852 DFRRQJI3VX1 $T=79520 87360 1 0 $X=79090 $Y=82240
X8735 1 2 241 346 84 110 DFRRQJI3VX1 $T=99680 150080 0 180 $X=84130 $Y=144960
X8736 1 2 241 358 84 840 DFRRQJI3VX1 $T=100240 150080 1 180 $X=84690 $Y=149440
X8737 1 2 241 359 84 1064 DFRRQJI3VX1 $T=100240 159040 0 180 $X=84690 $Y=153920
X8738 1 2 241 360 84 354 DFRRQJI3VX1 $T=85680 159040 0 0 $X=85250 $Y=158400
X8739 1 2 241 365 84 841 DFRRQJI3VX1 $T=100800 168000 0 180 $X=85250 $Y=162880
X8740 1 2 241 1367 84 335 DFRRQJI3VX1 $T=100800 176960 0 180 $X=85250 $Y=171840
X8741 1 2 241 117 84 303 DFRRQJI3VX1 $T=101360 168000 1 180 $X=85810 $Y=167360
X8742 1 2 241 351 94 331 DFRRQJI3VX1 $T=104720 114240 1 180 $X=89170 $Y=113600
X8743 1 2 241 352 94 106 DFRRQJI3VX1 $T=104720 123200 0 180 $X=89170 $Y=118080
X8744 1 2 129 1338 94 856 DFRRQJI3VX1 $T=109200 33600 0 180 $X=93650 $Y=28480
X8745 1 2 129 361 94 1188 DFRRQJI3VX1 $T=109200 33600 1 180 $X=93650 $Y=32960
X8746 1 2 129 1069 94 115 DFRRQJI3VX1 $T=109760 42560 0 180 $X=94210 $Y=37440
X8747 1 2 241 356 94 1074 DFRRQJI3VX1 $T=109760 51520 0 180 $X=94210 $Y=46400
X8748 1 2 241 120 94 276 DFRRQJI3VX1 $T=109760 78400 1 180 $X=94210 $Y=77760
X8749 1 2 241 363 94 286 DFRRQJI3VX1 $T=109760 87360 1 180 $X=94210 $Y=86720
X8750 1 2 241 370 94 341 DFRRQJI3VX1 $T=109760 96320 0 180 $X=94210 $Y=91200
X8751 1 2 241 371 94 111 DFRRQJI3VX1 $T=110320 96320 1 180 $X=94770 $Y=95680
X8752 1 2 241 857 94 848 DFRRQJI3VX1 $T=110320 114240 0 180 $X=94770 $Y=109120
X8753 1 2 246 1340 84 116 DFRRQJI3VX1 $T=110320 203840 0 180 $X=94770 $Y=198720
X8754 1 2 246 1339 84 369 DFRRQJI3VX1 $T=110320 212800 0 180 $X=94770 $Y=207680
X8755 1 2 246 860 84 1071 DFRRQJI3VX1 $T=110320 221760 0 180 $X=94770 $Y=216640
X8756 1 2 129 403 84 381 DFRRQJI3VX1 $T=108080 168000 1 0 $X=107650 $Y=162880
X8757 1 2 129 125 84 1078 DFRRQJI3VX1 $T=108080 168000 0 0 $X=107650 $Y=167360
X8758 1 2 129 398 84 378 DFRRQJI3VX1 $T=108080 176960 0 0 $X=107650 $Y=176320
X8759 1 2 246 1225 84 379 DFRRQJI3VX1 $T=108080 203840 0 0 $X=107650 $Y=203200
X8760 1 2 246 380 84 863 DFRRQJI3VX1 $T=108080 212800 0 0 $X=107650 $Y=212160
X8761 1 2 129 862 94 383 DFRRQJI3VX1 $T=109760 105280 1 0 $X=109330 $Y=100160
X8762 1 2 129 421 94 385 DFRRQJI3VX1 $T=110880 96320 1 0 $X=110450 $Y=91200
X8763 1 2 129 394 94 386 DFRRQJI3VX1 $T=110880 105280 0 0 $X=110450 $Y=104640
X8764 1 2 129 366 94 865 DFRRQJI3VX1 $T=111440 33600 1 0 $X=111010 $Y=28480
X8765 1 2 129 375 94 431 DFRRQJI3VX1 $T=111440 33600 0 0 $X=111010 $Y=32960
X8766 1 2 129 367 94 387 DFRRQJI3VX1 $T=111440 42560 1 0 $X=111010 $Y=37440
X8767 1 2 129 399 94 388 DFRRQJI3VX1 $T=111440 42560 0 0 $X=111010 $Y=41920
X8768 1 2 129 400 94 406 DFRRQJI3VX1 $T=111440 51520 0 0 $X=111010 $Y=50880
X8769 1 2 129 437 94 389 DFRRQJI3VX1 $T=111440 87360 0 0 $X=111010 $Y=86720
X8770 1 2 129 401 94 384 DFRRQJI3VX1 $T=112000 51520 1 0 $X=111570 $Y=46400
X8771 1 2 129 377 94 1016 DFRRQJI3VX1 $T=112560 114240 1 0 $X=112130 $Y=109120
X8772 1 2 129 395 84 864 DFRRQJI3VX1 $T=117600 185920 1 0 $X=117170 $Y=180800
X8773 1 2 129 408 84 128 DFRRQJI3VX1 $T=133280 176960 0 180 $X=117730 $Y=171840
X8774 1 2 246 418 84 426 DFRRQJI3VX1 $T=122640 221760 1 0 $X=122210 $Y=216640
X8775 1 2 129 448 84 433 DFRRQJI3VX1 $T=127120 168000 1 0 $X=126690 $Y=162880
X8776 1 2 129 397 84 1342 DFRRQJI3VX1 $T=127120 168000 0 0 $X=126690 $Y=167360
X8777 1 2 129 435 94 390 DFRRQJI3VX1 $T=143360 87360 1 180 $X=127810 $Y=86720
X8778 1 2 132 427 94 861 DFRRQJI3VX1 $T=143360 105280 0 180 $X=127810 $Y=100160
X8779 1 2 129 422 94 391 DFRRQJI3VX1 $T=143360 105280 1 180 $X=127810 $Y=104640
X8780 1 2 129 441 94 393 DFRRQJI3VX1 $T=143360 114240 0 180 $X=127810 $Y=109120
X8781 1 2 129 1098 94 413 DFRRQJI3VX1 $T=143920 42560 0 180 $X=128370 $Y=37440
X8782 1 2 129 415 94 446 DFRRQJI3VX1 $T=128800 42560 0 0 $X=128370 $Y=41920
X8783 1 2 129 443 94 442 DFRRQJI3VX1 $T=128800 51520 1 0 $X=128370 $Y=46400
X8784 1 2 129 416 94 1086 DFRRQJI3VX1 $T=128800 51520 0 0 $X=128370 $Y=50880
X8785 1 2 129 424 84 1067 DFRRQJI3VX1 $T=143920 123200 0 180 $X=128370 $Y=118080
X8786 1 2 129 449 84 409 DFRRQJI3VX1 $T=145040 176960 1 180 $X=129490 $Y=176320
X8787 1 2 129 417 94 459 DFRRQJI3VX1 $T=133280 60480 1 0 $X=132850 $Y=55360
X8788 1 2 129 432 94 429 DFRRQJI3VX1 $T=148400 60480 1 180 $X=132850 $Y=59840
X8789 1 2 132 411 94 438 DFRRQJI3VX1 $T=133280 69440 1 0 $X=132850 $Y=64320
X8790 1 2 129 439 84 404 DFRRQJI3VX1 $T=148400 159040 0 180 $X=132850 $Y=153920
X8791 1 2 246 1343 84 452 DFRRQJI3VX1 $T=138880 212800 0 0 $X=138450 $Y=212160
X8792 1 2 246 874 84 882 DFRRQJI3VX1 $T=138880 221760 1 0 $X=138450 $Y=216640
X8793 1 2 132 447 84 455 DFRRQJI3VX1 $T=139440 159040 0 0 $X=139010 $Y=158400
X8794 1 2 129 880 84 870 DFRRQJI3VX1 $T=155680 176960 0 180 $X=140130 $Y=171840
X8795 1 2 129 133 84 1085 DFRRQJI3VX1 $T=157360 168000 1 180 $X=141810 $Y=167360
X8796 1 2 132 463 84 423 DFRRQJI3VX1 $T=158480 105280 1 180 $X=142930 $Y=104640
X8797 1 2 132 1090 84 428 DFRRQJI3VX1 $T=159040 114240 1 180 $X=143490 $Y=113600
X8798 1 2 132 464 84 872 DFRRQJI3VX1 $T=159040 123200 0 180 $X=143490 $Y=118080
X8799 1 2 132 465 84 430 DFRRQJI3VX1 $T=159600 132160 1 180 $X=144050 $Y=131520
X8800 1 2 132 478 94 467 DFRRQJI3VX1 $T=145600 42560 1 0 $X=145170 $Y=37440
X8801 1 2 132 456 94 887 DFRRQJI3VX1 $T=145600 42560 0 0 $X=145170 $Y=41920
X8802 1 2 132 471 94 1346 DFRRQJI3VX1 $T=145600 51520 0 0 $X=145170 $Y=50880
X8803 1 2 132 468 84 436 DFRRQJI3VX1 $T=160720 150080 1 180 $X=145170 $Y=149440
X8804 1 2 132 475 94 1230 DFRRQJI3VX1 $T=163520 60480 0 180 $X=147970 $Y=55360
X8805 1 2 132 472 94 469 DFRRQJI3VX1 $T=163520 60480 1 180 $X=147970 $Y=59840
X8806 1 2 132 453 94 479 DFRRQJI3VX1 $T=148400 69440 1 0 $X=147970 $Y=64320
X8807 1 2 132 458 84 1234 DFRRQJI3VX1 $T=148400 159040 1 0 $X=147970 $Y=153920
X8808 1 2 246 1347 84 886 DFRRQJI3VX1 $T=170240 212800 1 180 $X=154690 $Y=212160
X8809 1 2 132 892 84 884 DFRRQJI3VX1 $T=170800 159040 1 180 $X=155250 $Y=158400
X8810 1 2 246 1096 84 482 DFRRQJI3VX1 $T=155680 212800 1 0 $X=155250 $Y=207680
X8811 1 2 129 1100 84 1093 DFRRQJI3VX1 $T=171360 176960 0 180 $X=155810 $Y=171840
X8812 1 2 129 1190 84 476 DFRRQJI3VX1 $T=171360 176960 1 180 $X=155810 $Y=176320
X8813 1 2 132 492 84 895 DFRRQJI3VX1 $T=156800 168000 1 0 $X=156370 $Y=162880
X8814 1 2 132 487 94 1097 DFRRQJI3VX1 $T=174160 33600 1 180 $X=158610 $Y=32960
X8815 1 2 132 894 94 481 DFRRQJI3VX1 $T=177520 42560 1 180 $X=161970 $Y=41920
X8816 1 2 147 486 94 899 DFRRQJI3VX1 $T=162960 51520 1 0 $X=162530 $Y=46400
X8817 1 2 132 144 94 137 DFRRQJI3VX1 $T=178080 51520 1 180 $X=162530 $Y=50880
X8818 1 2 132 504 94 1099 DFRRQJI3VX1 $T=178640 60480 0 180 $X=163090 $Y=55360
X8819 1 2 147 509 94 1237 DFRRQJI3VX1 $T=163520 60480 0 0 $X=163090 $Y=59840
X8820 1 2 147 508 94 491 DFRRQJI3VX1 $T=163520 69440 1 0 $X=163090 $Y=64320
X8821 1 2 132 510 94 140 DFRRQJI3VX1 $T=178640 69440 1 180 $X=163090 $Y=68800
X8822 1 2 246 499 184 496 DFRRQJI3VX1 $T=187040 212800 0 180 $X=171490 $Y=207680
X8823 1 2 246 1348 184 150 DFRRQJI3VX1 $T=171920 212800 0 0 $X=171490 $Y=212160
X8824 1 2 246 490 184 1108 DFRRQJI3VX1 $T=172480 203840 0 0 $X=172050 $Y=203200
X8825 1 2 132 149 184 483 DFRRQJI3VX1 $T=188160 159040 1 180 $X=172610 $Y=158400
X8826 1 2 132 503 184 484 DFRRQJI3VX1 $T=188160 168000 1 180 $X=172610 $Y=167360
X8827 1 2 132 513 184 1103 DFRRQJI3VX1 $T=188160 176960 0 180 $X=172610 $Y=171840
X8828 1 2 147 495 184 1109 DFRRQJI3VX1 $T=173040 176960 0 0 $X=172610 $Y=176320
X8829 1 2 246 516 184 493 DFRRQJI3VX1 $T=188160 185920 0 180 $X=172610 $Y=180800
X8830 1 2 147 905 94 900 DFRRQJI3VX1 $T=194320 42560 1 180 $X=178770 $Y=41920
X8831 1 2 147 143 94 994 DFRRQJI3VX1 $T=179200 69440 1 0 $X=178770 $Y=64320
X8832 1 2 147 521 94 511 DFRRQJI3VX1 $T=194880 51520 0 180 $X=179330 $Y=46400
X8833 1 2 147 522 94 507 DFRRQJI3VX1 $T=194880 51520 1 180 $X=179330 $Y=50880
X8834 1 2 147 1192 94 520 DFRRQJI3VX1 $T=179760 60480 0 0 $X=179330 $Y=59840
X8835 1 2 147 517 94 1307 DFRRQJI3VX1 $T=179760 69440 0 0 $X=179330 $Y=68800
X8836 1 2 147 632 94 494 DFRRQJI3VX1 $T=197680 114240 0 180 $X=182130 $Y=109120
X8837 1 2 147 571 94 497 DFRRQJI3VX1 $T=197680 114240 1 180 $X=182130 $Y=113600
X8838 1 2 147 606 94 1106 DFRRQJI3VX1 $T=197680 123200 1 180 $X=182130 $Y=122560
X8839 1 2 147 586 184 498 DFRRQJI3VX1 $T=197680 132160 1 180 $X=182130 $Y=131520
X8840 1 2 147 552 184 134 DFRRQJI3VX1 $T=197680 141120 1 180 $X=182130 $Y=140480
X8841 1 2 246 529 184 528 DFRRQJI3VX1 $T=188160 212800 1 0 $X=187730 $Y=207680
X8842 1 2 246 1370 184 527 DFRRQJI3VX1 $T=188720 203840 0 0 $X=188290 $Y=203200
X8843 1 2 147 530 184 515 DFRRQJI3VX1 $T=204960 185920 0 180 $X=189410 $Y=180800
X8844 1 2 147 535 184 911 DFRRQJI3VX1 $T=190960 150080 1 0 $X=190530 $Y=144960
X8845 1 2 147 578 184 901 DFRRQJI3VX1 $T=206080 168000 0 180 $X=190530 $Y=162880
X8846 1 2 147 579 184 155 DFRRQJI3VX1 $T=206080 168000 1 180 $X=190530 $Y=167360
X8847 1 2 147 156 184 902 DFRRQJI3VX1 $T=206080 176960 0 180 $X=190530 $Y=171840
X8848 1 2 147 551 184 500 DFRRQJI3VX1 $T=206640 141120 0 180 $X=191090 $Y=136000
X8849 1 2 147 512 184 525 DFRRQJI3VX1 $T=206640 159040 1 180 $X=191090 $Y=158400
X8850 1 2 147 907 184 995 DFRRQJI3VX1 $T=191520 176960 0 0 $X=191090 $Y=176320
X8851 1 2 147 533 94 523 DFRRQJI3VX1 $T=211120 69440 0 180 $X=195570 $Y=64320
X8852 1 2 147 160 94 1308 DFRRQJI3VX1 $T=211120 78400 0 180 $X=195570 $Y=73280
X8853 1 2 147 158 94 1309 DFRRQJI3VX1 $T=211680 42560 1 180 $X=196130 $Y=41920
X8854 1 2 147 1311 94 910 DFRRQJI3VX1 $T=211680 51520 0 180 $X=196130 $Y=46400
X8855 1 2 147 1193 94 543 DFRRQJI3VX1 $T=211680 51520 1 180 $X=196130 $Y=50880
X8856 1 2 147 1110 94 904 DFRRQJI3VX1 $T=211680 60480 0 180 $X=196130 $Y=55360
X8857 1 2 147 1363 94 903 DFRRQJI3VX1 $T=211680 69440 1 180 $X=196130 $Y=68800
X8858 1 2 147 157 94 539 DFRRQJI3VX1 $T=211680 78400 1 180 $X=196130 $Y=77760
X8859 1 2 147 580 94 519 DFRRQJI3VX1 $T=212240 105280 0 180 $X=196690 $Y=100160
X8860 1 2 147 581 94 524 DFRRQJI3VX1 $T=213920 114240 0 180 $X=198370 $Y=109120
X8861 1 2 147 576 94 526 DFRRQJI3VX1 $T=213920 114240 1 180 $X=198370 $Y=113600
X8862 1 2 246 913 184 1113 DFRRQJI3VX1 $T=215040 212800 1 180 $X=199490 $Y=212160
X8863 1 2 568 555 178 174 DFRRQJI3VX1 $T=213920 51520 0 0 $X=213490 $Y=50880
X8864 1 2 568 161 184 165 DFRRQJI3VX1 $T=213920 168000 1 0 $X=213490 $Y=162880
X8865 1 2 147 162 184 559 DFRRQJI3VX1 $T=213920 168000 0 0 $X=213490 $Y=167360
X8866 1 2 568 1194 184 171 DFRRQJI3VX1 $T=213920 176960 1 0 $X=213490 $Y=171840
X8867 1 2 181 573 184 544 DFRRQJI3VX1 $T=213920 185920 1 0 $X=213490 $Y=180800
X8868 1 2 181 1349 184 915 DFRRQJI3VX1 $T=213920 212800 1 0 $X=213490 $Y=207680
X8869 1 2 568 569 178 560 DFRRQJI3VX1 $T=214480 42560 0 0 $X=214050 $Y=41920
X8870 1 2 568 163 178 1120 DFRRQJI3VX1 $T=214480 51520 1 0 $X=214050 $Y=46400
X8871 1 2 568 164 178 561 DFRRQJI3VX1 $T=214480 60480 1 0 $X=214050 $Y=55360
X8872 1 2 568 166 178 917 DFRRQJI3VX1 $T=214480 60480 0 0 $X=214050 $Y=59840
X8873 1 2 568 169 178 1245 DFRRQJI3VX1 $T=214480 69440 1 0 $X=214050 $Y=64320
X8874 1 2 568 575 178 562 DFRRQJI3VX1 $T=214480 69440 0 0 $X=214050 $Y=68800
X8875 1 2 568 574 178 563 DFRRQJI3VX1 $T=214480 78400 1 0 $X=214050 $Y=73280
X8876 1 2 568 168 178 1244 DFRRQJI3VX1 $T=214480 78400 0 0 $X=214050 $Y=77760
X8877 1 2 181 916 184 557 DFRRQJI3VX1 $T=217840 212800 0 0 $X=217410 $Y=212160
X8878 1 2 181 597 184 1196 DFRRQJI3VX1 $T=226800 176960 0 0 $X=226370 $Y=176320
X8879 1 2 181 923 184 587 DFRRQJI3VX1 $T=244160 168000 1 180 $X=228610 $Y=167360
X8880 1 2 181 595 184 1129 DFRRQJI3VX1 $T=229040 176960 1 0 $X=228610 $Y=171840
X8881 1 2 181 585 184 570 DFRRQJI3VX1 $T=246400 212800 0 180 $X=230850 $Y=207680
X8882 1 2 568 611 178 1250 DFRRQJI3VX1 $T=231840 78400 1 0 $X=231410 $Y=73280
X8883 1 2 568 627 178 601 DFRRQJI3VX1 $T=231840 78400 0 0 $X=231410 $Y=77760
X8884 1 2 568 590 178 1126 DFRRQJI3VX1 $T=247520 42560 1 180 $X=231970 $Y=41920
X8885 1 2 568 605 178 919 DFRRQJI3VX1 $T=247520 51520 0 180 $X=231970 $Y=46400
X8886 1 2 568 600 178 589 DFRRQJI3VX1 $T=232400 51520 0 0 $X=231970 $Y=50880
X8887 1 2 568 189 178 1125 DFRRQJI3VX1 $T=247520 60480 0 180 $X=231970 $Y=55360
X8888 1 2 568 179 178 926 DFRRQJI3VX1 $T=232960 60480 0 0 $X=232530 $Y=59840
X8889 1 2 568 610 178 1124 DFRRQJI3VX1 $T=248080 69440 0 180 $X=232530 $Y=64320
X8890 1 2 568 175 178 593 DFRRQJI3VX1 $T=248080 69440 1 180 $X=232530 $Y=68800
X8891 1 2 181 592 184 572 DFRRQJI3VX1 $T=253680 194880 1 180 $X=238130 $Y=194240
X8892 1 2 181 604 184 588 DFRRQJI3VX1 $T=253680 203840 1 180 $X=238130 $Y=203200
X8893 1 2 181 997 184 172 DFRRQJI3VX1 $T=255920 185920 0 180 $X=240370 $Y=180800
X8894 1 2 181 183 184 1253 DFRRQJI3VX1 $T=241360 185920 0 0 $X=240930 $Y=185280
X8895 1 2 181 187 184 924 DFRRQJI3VX1 $T=257040 176960 1 180 $X=241490 $Y=176320
X8896 1 2 568 191 178 927 DFRRQJI3VX1 $T=265440 51520 0 180 $X=249890 $Y=46400
X8897 1 2 568 618 178 928 DFRRQJI3VX1 $T=265440 51520 1 180 $X=249890 $Y=50880
X8898 1 2 568 626 178 186 DFRRQJI3VX1 $T=265440 60480 0 180 $X=249890 $Y=55360
X8899 1 2 568 625 178 1356 DFRRQJI3VX1 $T=250320 69440 1 0 $X=249890 $Y=64320
X8900 1 2 568 628 178 1254 DFRRQJI3VX1 $T=250320 69440 0 0 $X=249890 $Y=68800
X8901 1 2 568 614 178 599 DFRRQJI3VX1 $T=267120 105280 0 180 $X=251570 $Y=100160
X8902 1 2 181 631 184 598 DFRRQJI3VX1 $T=273280 185920 1 180 $X=257730 $Y=185280
X8903 1 2 643 615 184 933 DFRRQJI3VX1 $T=258720 185920 1 0 $X=258290 $Y=180800
X8904 1 2 657 1140 188 1146 DFRRQJI3VX1 $T=266000 203840 0 0 $X=265570 $Y=203200
X8905 1 2 657 1256 188 642 DFRRQJI3VX1 $T=266000 212800 0 0 $X=265570 $Y=212160
X8906 1 2 181 193 178 939 DFRRQJI3VX1 $T=267120 105280 1 0 $X=266690 $Y=100160
X8907 1 2 568 935 178 636 DFRRQJI3VX1 $T=282800 51520 0 180 $X=267250 $Y=46400
X8908 1 2 568 645 178 932 DFRRQJI3VX1 $T=282800 51520 1 180 $X=267250 $Y=50880
X8909 1 2 568 654 178 937 DFRRQJI3VX1 $T=267680 60480 1 0 $X=267250 $Y=55360
X8910 1 2 568 665 178 623 DFRRQJI3VX1 $T=282800 60480 1 180 $X=267250 $Y=59840
X8911 1 2 568 652 178 194 DFRRQJI3VX1 $T=282800 69440 0 180 $X=267250 $Y=64320
X8912 1 2 568 658 178 629 DFRRQJI3VX1 $T=282800 69440 1 180 $X=267250 $Y=68800
X8913 1 2 568 635 178 1260 DFRRQJI3VX1 $T=269360 42560 1 0 $X=268930 $Y=37440
X8914 1 2 219 660 178 649 DFRRQJI3VX1 $T=272160 78400 1 0 $X=271730 $Y=73280
X8915 1 2 219 704 178 653 DFRRQJI3VX1 $T=292320 114240 1 180 $X=276770 $Y=113600
X8916 1 2 657 1147 188 663 DFRRQJI3VX1 $T=277200 194880 0 0 $X=276770 $Y=194240
X8917 1 2 672 941 184 1155 DFRRQJI3VX1 $T=279440 185920 1 0 $X=279010 $Y=180800
X8918 1 2 938 675 184 1259 DFRRQJI3VX1 $T=295120 176960 0 180 $X=279570 $Y=171840
X8919 1 2 657 673 188 669 DFRRQJI3VX1 $T=297920 203840 1 180 $X=282370 $Y=203200
X8920 1 2 1263 667 184 1156 DFRRQJI3VX1 $T=283920 168000 0 0 $X=283490 $Y=167360
X8921 1 2 657 1357 188 656 DFRRQJI3VX1 $T=299040 212800 1 180 $X=283490 $Y=212160
X8922 1 2 650 677 184 655 DFRRQJI3VX1 $T=299600 168000 0 180 $X=284050 $Y=162880
X8923 1 2 672 1150 184 942 DFRRQJI3VX1 $T=284480 185920 0 0 $X=284050 $Y=185280
X8924 1 2 568 684 178 1149 DFRRQJI3VX1 $T=300160 42560 1 180 $X=284610 $Y=41920
X8925 1 2 568 201 178 668 DFRRQJI3VX1 $T=300160 51520 0 180 $X=284610 $Y=46400
X8926 1 2 568 678 178 940 DFRRQJI3VX1 $T=300160 51520 1 180 $X=284610 $Y=50880
X8927 1 2 219 689 178 1323 DFRRQJI3VX1 $T=285040 60480 1 0 $X=284610 $Y=55360
X8928 1 2 219 694 178 1266 DFRRQJI3VX1 $T=285040 69440 1 0 $X=284610 $Y=64320
X8929 1 2 219 661 178 679 DFRRQJI3VX1 $T=285040 69440 0 0 $X=284610 $Y=68800
X8930 1 2 219 690 178 948 DFRRQJI3VX1 $T=294000 96320 0 0 $X=293570 $Y=95680
X8931 1 2 219 691 178 1270 DFRRQJI3VX1 $T=294000 105280 1 0 $X=293570 $Y=100160
X8932 1 2 219 707 178 676 DFRRQJI3VX1 $T=309680 87360 0 180 $X=294130 $Y=82240
X8933 1 2 219 695 178 1152 DFRRQJI3VX1 $T=309680 96320 0 180 $X=294130 $Y=91200
X8934 1 2 712 1157 184 1411 DFRRQJI3VX1 $T=297920 203840 1 0 $X=297490 $Y=198720
X8935 1 2 943 1358 184 700 DFRRQJI3VX1 $T=313600 203840 1 180 $X=298050 $Y=203200
X8936 1 2 949 203 184 685 DFRRQJI3VX1 $T=315840 159040 1 180 $X=300290 $Y=158400
X8937 1 2 1160 702 184 1161 DFRRQJI3VX1 $T=300720 168000 1 0 $X=300290 $Y=162880
X8938 1 2 219 1359 178 1158 DFRRQJI3VX1 $T=316960 51520 0 180 $X=301410 $Y=46400
X8939 1 2 219 1199 178 945 DFRRQJI3VX1 $T=316960 51520 1 180 $X=301410 $Y=50880
X8940 1 2 219 741 178 710 DFRRQJI3VX1 $T=316960 60480 1 180 $X=301410 $Y=59840
X8941 1 2 219 740 178 693 DFRRQJI3VX1 $T=316960 69440 0 180 $X=301410 $Y=64320
X8942 1 2 219 952 184 946 DFRRQJI3VX1 $T=317520 159040 0 180 $X=301970 $Y=153920
X8943 1 2 697 714 184 209 DFRRQJI3VX1 $T=322000 212800 0 180 $X=306450 $Y=207680
X8944 1 2 1269 210 184 703 DFRRQJI3VX1 $T=322000 212800 1 180 $X=306450 $Y=212160
X8945 1 2 219 729 178 222 DFRRQJI3VX1 $T=319760 51520 0 0 $X=319330 $Y=50880
X8946 1 2 219 1174 178 725 DFRRQJI3VX1 $T=319760 60480 1 0 $X=319330 $Y=55360
X8947 1 2 219 213 178 1275 DFRRQJI3VX1 $T=319760 60480 0 0 $X=319330 $Y=59840
X8948 1 2 219 742 178 1167 DFRRQJI3VX1 $T=319760 69440 1 0 $X=319330 $Y=64320
X8949 1 2 219 211 178 727 DFRRQJI3VX1 $T=319760 96320 1 0 $X=319330 $Y=91200
X8950 1 2 219 216 178 1163 DFRRQJI3VX1 $T=319760 96320 0 0 $X=319330 $Y=95680
X8951 1 2 219 718 178 726 DFRRQJI3VX1 $T=319760 105280 1 0 $X=319330 $Y=100160
X8952 1 2 219 716 178 728 DFRRQJI3VX1 $T=319760 114240 1 0 $X=319330 $Y=109120
X8953 1 2 219 743 184 207 DFRRQJI3VX1 $T=319760 141120 1 0 $X=319330 $Y=136000
X8954 1 2 219 214 184 208 DFRRQJI3VX1 $T=319760 141120 0 0 $X=319330 $Y=140480
X8955 1 2 219 1200 184 217 DFRRQJI3VX1 $T=319760 150080 0 0 $X=319330 $Y=149440
X8956 1 2 226 720 184 1380 DFRRQJI3VX1 $T=319760 159040 0 0 $X=319330 $Y=158400
X8957 1 2 733 737 184 961 DFRRQJI3VX1 $T=319760 168000 1 0 $X=319330 $Y=162880
X8958 1 2 226 752 184 1329 DFRRQJI3VX1 $T=334880 141120 0 0 $X=334450 $Y=140480
X8959 1 2 226 980 184 1276 DFRRQJI3VX1 $T=350000 150080 1 180 $X=334450 $Y=149440
X8960 1 2 219 753 178 1171 DFRRQJI3VX1 $T=351680 42560 1 180 $X=336130 $Y=41920
X8961 1 2 219 754 178 962 DFRRQJI3VX1 $T=351680 51520 0 180 $X=336130 $Y=46400
X8962 1 2 219 1328 178 1279 DFRRQJI3VX1 $T=351680 51520 1 180 $X=336130 $Y=50880
X8963 1 2 219 756 178 223 DFRRQJI3VX1 $T=351680 60480 1 180 $X=336130 $Y=59840
X8964 1 2 219 751 178 1288 DFRRQJI3VX1 $T=336560 105280 1 0 $X=336130 $Y=100160
X8965 1 2 219 747 178 968 DFRRQJI3VX1 $T=352240 69440 0 180 $X=336690 $Y=64320
X8966 1 2 219 739 178 1287 DFRRQJI3VX1 $T=337120 96320 0 0 $X=336690 $Y=95680
X8967 1 2 219 759 178 1327 DFRRQJI3VX1 $T=360080 69440 1 180 $X=344530 $Y=68800
X8968 1 2 219 755 178 1282 DFRRQJI3VX1 $T=360080 78400 0 180 $X=344530 $Y=73280
X8969 1 2 219 1182 178 762 DFRRQJI3VX1 $T=344960 87360 0 0 $X=344530 $Y=86720
X8970 1 2 226 764 184 744 DFRRQJI3VX1 $T=361200 159040 1 180 $X=345650 $Y=158400
X8971 1 2 226 1201 184 745 DFRRQJI3VX1 $T=361200 168000 0 180 $X=345650 $Y=162880
X8972 1 2 226 748 184 984 DFRRQJI3VX1 $T=346640 150080 1 0 $X=346210 $Y=144960
X8973 1 2 226 231 184 763 DFRRQJI3VX1 $T=346640 159040 1 0 $X=346210 $Y=153920
X8974 1 2 226 769 184 974 DFRRQJI3VX1 $T=361760 168000 1 180 $X=346210 $Y=167360
X8975 1 2 219 234 178 982 DFRRQJI3VX1 $T=367360 60480 1 180 $X=351810 $Y=59840
X8976 1 2 219 757 178 1331 DFRRQJI3VX1 $T=352240 69440 1 0 $X=351810 $Y=64320
X8977 1 2 1289 1203 184 758 DFRRQJI3VX1 $T=367360 203840 0 180 $X=351810 $Y=198720
X8978 1 2 219 777 178 225 DFRRQJI3VX1 $T=367920 51520 1 180 $X=352370 $Y=50880
X8979 1 2 983 1202 184 1179 DFRRQJI3VX1 $T=371280 194880 1 180 $X=355730 $Y=194240
X8980 1 2 226 233 178 1293 DFRRQJI3VX1 $T=363440 78400 1 0 $X=363010 $Y=73280
X8981 1 2 226 232 178 772 DFRRQJI3VX1 $T=378560 78400 1 180 $X=363010 $Y=77760
X8982 1 2 226 770 178 1295 DFRRQJI3VX1 $T=363440 87360 0 0 $X=363010 $Y=86720
X8983 1 2 226 784 178 986 DFRRQJI3VX1 $T=363440 96320 1 0 $X=363010 $Y=91200
X8984 1 2 226 786 184 765 DFRRQJI3VX1 $T=378560 150080 1 180 $X=363010 $Y=149440
X8985 1 2 226 785 184 1294 DFRRQJI3VX1 $T=363440 159040 1 0 $X=363010 $Y=153920
X8986 1 2 219 787 178 229 DFRRQJI3VX1 $T=379120 42560 0 180 $X=363570 $Y=37440
X8987 1 2 219 788 178 1290 DFRRQJI3VX1 $T=379120 42560 1 180 $X=363570 $Y=41920
X8988 1 2 219 778 178 228 DFRRQJI3VX1 $T=379120 51520 0 180 $X=363570 $Y=46400
X8989 1 2 219 779 178 761 DFRRQJI3VX1 $T=379120 60480 0 180 $X=363570 $Y=55360
X8990 1 2 219 782 178 985 DFRRQJI3VX1 $T=364000 69440 0 0 $X=363570 $Y=68800
X8991 1 2 226 775 184 1184 DFRRQJI3VX1 $T=364000 159040 0 0 $X=363570 $Y=158400
X8992 1 2 226 789 184 1181 DFRRQJI3VX1 $T=379120 168000 0 180 $X=363570 $Y=162880
X8993 1 2 226 780 184 1180 DFRRQJI3VX1 $T=379120 168000 1 180 $X=363570 $Y=167360
X8994 1 2 219 781 178 1412 DFRRQJI3VX1 $T=379680 33600 1 180 $X=364130 $Y=32960
X8995 1 2 219 783 178 236 DFRRQJI3VX1 $T=367360 69440 1 0 $X=366930 $Y=64320
X8996 1 2 802 1413 1210 271 987 ON211JI3VX1 $T=53200 69440 0 180 $X=48850 $Y=64320
X8997 1 2 96 1213 804 270 283 ON211JI3VX1 $T=52080 51520 0 0 $X=51650 $Y=50880
X8998 1 2 283 1027 87 271 enable ON211JI3VX1 $T=54320 60480 0 0 $X=53890 $Y=59840
X8999 1 2 303 1029 1033 1028 811 ON211JI3VX1 $T=58800 185920 0 180 $X=54450 $Y=180800
X9000 1 2 113 1030 1392 814 810 ON211JI3VX1 $T=60480 96320 0 180 $X=56130 $Y=91200
X9001 1 2 113 99 1366 818 1036 ON211JI3VX1 $T=65520 96320 0 180 $X=61170 $Y=91200
X9002 1 2 297 1301 1414 820 300 ON211JI3VX1 $T=62160 185920 1 0 $X=61730 $Y=180800
X9003 1 2 113 1042 294 822 821 ON211JI3VX1 $T=71120 96320 0 180 $X=66770 $Y=91200
X9004 1 2 303 1220 1053 311 1050 ON211JI3VX1 $T=75040 185920 0 0 $X=74610 $Y=185280
X9005 1 2 1057 340 1415 320 837 ON211JI3VX1 $T=80080 176960 0 0 $X=79650 $Y=176320
X9006 1 2 enable 1416 372 853 113 ON211JI3VX1 $T=105280 176960 1 180 $X=100930 $Y=176320
X9007 1 2 460 1375 1087 466 1304 ON211JI3VX1 $T=151200 185920 1 180 $X=146850 $Y=185280
X9008 1 2 995 1312 1417 538 906 ON211JI3VX1 $T=204400 194880 1 180 $X=200050 $Y=194240
X9009 1 2 1156 205 696 947 200 ON211JI3VX1 $T=301840 176960 1 0 $X=301410 $Y=171840
X9010 1 2 749 963 1391 1325 730 ON211JI3VX1 $T=331520 176960 1 0 $X=331090 $Y=171840
X9011 1 2 218 723 1169 960 enable ON211JI3VX1 $T=335440 185920 0 180 $X=331090 $Y=180800
X9012 1 2 1012 87 1006 86 247 ON22JI3VX1 $T=34720 69440 1 180 $X=29810 $Y=68800
X9013 1 2 131 98 1186 807 305 ON22JI3VX1 $T=57120 42560 0 180 $X=52210 $Y=37440
X9014 1 2 293 1043 1418 833 1037 ON22JI3VX1 $T=69440 203840 1 180 $X=64530 $Y=203200
X9015 1 2 1085 414 1419 876 870 ON22JI3VX1 $T=140560 185920 1 0 $X=140130 $Y=180800
X9016 1 2 878 136 1343 877 876 ON22JI3VX1 $T=148960 203840 1 180 $X=144050 $Y=203200
X9017 1 2 885 136 1347 1344 1094 ON22JI3VX1 $T=156800 203840 0 0 $X=156370 $Y=203200
X9018 1 2 993 136 1348 898 1104 ON22JI3VX1 $T=179760 203840 0 180 $X=174850 $Y=198720
X9019 1 2 527 167 1370 541 152 ON22JI3VX1 $T=189280 203840 1 0 $X=188850 $Y=198720
X9020 1 2 527 1239 537 152 528 ON22JI3VX1 $T=193760 203840 1 0 $X=193330 $Y=198720
X9021 1 2 915 556 1350 173 557 ON22JI3VX1 $T=220080 194880 0 0 $X=219650 $Y=194240
X9022 1 2 570 1122 585 920 176 ON22JI3VX1 $T=229600 203840 0 0 $X=229170 $Y=203200
X9023 1 2 598 1420 922 925 924 ON22JI3VX1 $T=246400 194880 0 180 $X=241490 $Y=189760
X9024 1 2 1153 1154 1358 713 950 ON22JI3VX1 $T=304640 194880 1 0 $X=304210 $Y=189760
X9025 1 2 209 206 955 732 703 ON22JI3VX1 $T=316960 185920 1 180 $X=312050 $Y=185280
X9026 1 2 961 958 1165 722 217 ON22JI3VX1 $T=324800 185920 1 0 $X=324370 $Y=180800
X9027 1 2 758 738 1373 970 1179 ON22JI3VX1 $T=347200 194880 1 0 $X=346770 $Y=189760
X9028 1 2 1181 1001 760 1330 1180 ON22JI3VX1 $T=361200 176960 0 180 $X=356290 $Y=171840
X9029 1 2 226 1292 184 981 DFRRQJI3VX2 $T=372400 194880 0 180 $X=355730 $Y=189760
X9030 1 2 386 88 253 244 EO3JI3VX1 $T=49840 105280 0 180 $X=38770 $Y=100160
X9031 1 2 386 91 1207 1185 EO3JI3VX1 $T=53760 105280 1 180 $X=42690 $Y=104640
X9032 1 2 1015 796 98 NO2JI3VX0 $T=44800 51520 0 180 $X=42130 $Y=46400
X9033 1 2 1421 1015 1027 NO2JI3VX0 $T=43120 60480 0 0 $X=42690 $Y=59840
X9034 1 2 798 255 257 NO2JI3VX0 $T=43120 78400 1 0 $X=42690 $Y=73280
X9035 1 2 807 1023 90 NO2JI3VX0 $T=52640 42560 0 180 $X=49970 $Y=37440
X9036 1 2 1422 1210 96 NO2JI3VX0 $T=51520 60480 1 0 $X=51090 $Y=55360
X9037 1 2 260 988 322 NO2JI3VX0 $T=51520 203840 1 0 $X=51090 $Y=198720
X9038 1 2 808 807 98 NO2JI3VX0 $T=52640 42560 0 0 $X=52210 $Y=41920
X9039 1 2 279 1033 1034 NO2JI3VX0 $T=61040 176960 1 180 $X=58370 $Y=176320
X9040 1 2 292 1187 1045 NO2JI3VX0 $T=68320 194880 1 0 $X=67890 $Y=189760
X9041 1 2 826 1415 297 NO2JI3VX0 $T=71680 176960 0 0 $X=71250 $Y=176320
X9042 1 2 830 105 267 NO2JI3VX0 $T=76720 212800 0 180 $X=74050 $Y=207680
X9043 1 2 347 830 308 NO2JI3VX0 $T=80080 212800 0 180 $X=77410 $Y=207680
X9044 1 2 1070 345 848 NO2JI3VX0 $T=95200 114240 0 180 $X=92530 $Y=109120
X9045 1 2 124 127 126 NO2JI3VX0 $T=113120 194880 1 0 $X=112690 $Y=189760
X9046 1 2 369 1368 116 NO2JI3VX0 $T=113120 194880 0 0 $X=112690 $Y=194240
X9047 1 2 307 505 126 NO2JI3VX0 $T=131600 194880 1 180 $X=128930 $Y=194240
X9048 1 2 1231 445 451 NO2JI3VX0 $T=151760 194880 1 180 $X=149090 $Y=194240
X9049 1 2 451 881 884 NO2JI3VX0 $T=150640 194880 1 0 $X=150210 $Y=189760
X9050 1 2 1094 444 1093 NO2JI3VX0 $T=160720 185920 0 180 $X=158050 $Y=180800
X9051 1 2 139 135 477 NO2JI3VX0 $T=164080 194880 1 180 $X=161410 $Y=194240
X9052 1 2 502 896 1103 NO2JI3VX0 $T=175840 185920 1 180 $X=173170 $Y=185280
X9053 1 2 502 506 150 NO2JI3VX0 $T=185920 203840 0 180 $X=183250 $Y=198720
X9054 1 2 908 1314 559 NO2JI3VX0 $T=210560 194880 0 180 $X=207890 $Y=189760
X9055 1 2 556 1241 172 NO2JI3VX0 $T=224560 194880 0 0 $X=224130 $Y=194240
X9056 1 2 612 1423 1130 NO2JI3VX0 $T=246400 24640 0 0 $X=245970 $Y=24000
X9057 1 2 1251 1133 996 NO2JI3VX0 $T=250880 24640 0 0 $X=250450 $Y=24000
X9058 1 2 617 1135 609 NO2JI3VX0 $T=260960 33600 0 180 $X=258290 $Y=28480
X9059 1 2 177 1424 613 NO2JI3VX0 $T=263200 24640 1 180 $X=260530 $Y=24000
X9060 1 2 659 666 1148 NO2JI3VX0 $T=283360 212800 1 0 $X=282930 $Y=207680
X9061 1 2 1322 1357 666 NO2JI3VX0 $T=291760 212800 1 0 $X=291330 $Y=207680
X9062 1 2 1151 1154 126 NO2JI3VX0 $T=297360 194880 0 0 $X=296930 $Y=194240
X9063 1 2 713 1151 942 NO2JI3VX0 $T=302960 194880 1 180 $X=300290 $Y=194240
X9064 1 2 202 1159 946 NO2JI3VX0 $T=309680 185920 0 180 $X=307010 $Y=180800
X9065 1 2 696 705 202 NO2JI3VX0 $T=310800 185920 1 180 $X=308130 $Y=185280
X9066 1 2 954 1425 205 NO2JI3VX0 $T=313600 176960 0 0 $X=313170 $Y=176320
X9067 1 2 732 1175 206 NO2JI3VX0 $T=335440 185920 1 0 $X=335010 $Y=180800
X9068 1 2 1172 1170 744 NO2JI3VX0 $T=337680 185920 1 180 $X=335010 $Y=185280
X9069 1 2 206 227 1276 NO2JI3VX0 $T=338800 168000 1 180 $X=336130 $Y=167360
X9070 1 2 738 724 745 NO2JI3VX0 $T=343280 185920 0 180 $X=340610 $Y=180800
X9071 1 2 973 969 974 NO2JI3VX0 $T=347760 176960 0 180 $X=345090 $Y=171840
X9072 1 2 1408 86 1004 1011 ON21JI3VX1 $T=34720 60480 0 0 $X=34290 $Y=59840
X9073 1 2 247 255 1013 1012 ON21JI3VX1 $T=35840 69440 0 0 $X=35410 $Y=68800
X9074 1 2 1386 261 1007 1010 ON21JI3VX1 $T=40320 203840 1 180 $X=36530 $Y=203200
X9075 1 2 1009 255 794 1205 ON21JI3VX1 $T=44800 69440 0 180 $X=41010 $Y=64320
X9076 1 2 1409 274 1206 1020 ON21JI3VX1 $T=46480 33600 1 180 $X=42690 $Y=32960
X9077 1 2 1023 1186 1020 93 ON21JI3VX1 $T=51520 33600 1 180 $X=47730 $Y=32960
X9078 1 2 279 269 811 1034 ON21JI3VX1 $T=54320 176960 0 0 $X=53890 $Y=176320
X9079 1 2 988 1212 816 1299 ON21JI3VX1 $T=54320 194880 0 0 $X=53890 $Y=194240
X9080 1 2 305 274 819 1362 ON21JI3VX1 $T=61600 33600 0 0 $X=61170 $Y=32960
X9081 1 2 826 105 1048 989 ON21JI3VX1 $T=70560 203840 1 0 $X=70130 $Y=198720
X9082 1 2 1387 347 860 1337 ON21JI3VX1 $T=100240 212800 0 0 $X=99810 $Y=212160
X9083 1 2 180 1076 630 1374 ON21JI3VX1 $T=101920 24640 1 0 $X=101490 $Y=19520
X9084 1 2 859 355 1340 858 ON21JI3VX1 $T=105280 194880 1 180 $X=101490 $Y=194240
X9085 1 2 374 373 1341 372 ON21JI3VX1 $T=122080 185920 1 180 $X=118290 $Y=185280
X9086 1 2 1388 136 1081 1082 ON21JI3VX1 $T=132160 203840 1 180 $X=128370 $Y=203200
X9087 1 2 180 1426 934 1228 ON21JI3VX1 $T=129920 24640 0 0 $X=129490 $Y=24000
X9088 1 2 180 1427 651 871 ON21JI3VX1 $T=141120 33600 1 0 $X=140690 $Y=28480
X9089 1 2 180 1428 641 457 ON21JI3VX1 $T=154000 33600 0 0 $X=153570 $Y=32960
X9090 1 2 470 896 1429 480 ON21JI3VX1 $T=171920 194880 0 180 $X=168130 $Y=189760
X9091 1 2 502 898 490 1236 ON21JI3VX1 $T=171360 203840 1 0 $X=170930 $Y=198720
X9092 1 2 902 152 1238 531 ON21JI3VX1 $T=194320 194880 1 0 $X=193890 $Y=189760
X9093 1 2 180 1114 609 909 ON21JI3VX1 $T=201040 33600 1 0 $X=200610 $Y=28480
X9094 1 2 536 1389 1351 545 ON21JI3VX1 $T=207760 185920 0 0 $X=207330 $Y=185280
X9095 1 2 180 1430 613 1315 ON21JI3VX1 $T=221760 24640 0 0 $X=221330 $Y=24000
X9096 1 2 180 918 617 1243 ON21JI3VX1 $T=226240 33600 1 0 $X=225810 $Y=28480
X9097 1 2 566 1390 1195 1353 ON21JI3VX1 $T=227360 194880 1 0 $X=226930 $Y=189760
X9098 1 2 570 167 1248 920 ON21JI3VX1 $T=229600 203840 1 0 $X=229170 $Y=198720
X9099 1 2 180 1127 177 1247 ON21JI3VX1 $T=236320 33600 0 0 $X=235890 $Y=32960
X9100 1 2 180 1431 1251 1354 ON21JI3VX1 $T=239120 24640 1 0 $X=238690 $Y=19520
X9101 1 2 159 1248 1432 1316 ON21JI3VX1 $T=240800 203840 1 0 $X=240370 $Y=198720
X9102 1 2 180 1433 1130 1355 ON21JI3VX1 $T=247520 42560 0 180 $X=243730 $Y=37440
X9103 1 2 180 1318 996 1317 ON21JI3VX1 $T=256480 33600 1 180 $X=252690 $Y=32960
X9104 1 2 180 1136 612 1138 ON21JI3VX1 $T=258160 33600 0 0 $X=257730 $Y=32960
X9105 1 2 202 1154 1157 1268 ON21JI3VX1 $T=308000 194880 1 180 $X=304210 $Y=194240
X9106 1 2 1159 711 1377 692 ON21JI3VX1 $T=311360 176960 1 180 $X=307570 $Y=176320
X9107 1 2 713 1272 1277 1273 ON21JI3VX1 $T=329280 203840 0 0 $X=328850 $Y=203200
X9108 1 2 651 1095 1434 671 641 OR4JI3VX1 $T=286160 24640 1 180 $X=279570 $Y=24000
X9109 1 2 215 204 1271 701 688 OR4JI3VX1 $T=315840 33600 0 180 $X=309250 $Y=28480
X9110 1 2 736 1166 698 715 532 OR4JI3VX1 $T=331520 24640 1 180 $X=324930 $Y=24000
X9111 1 2 750 977 978 767 976 OR4JI3VX1 $T=353360 33600 0 180 $X=346770 $Y=28480
X9112 1 2 534 546 BUJI3VX16 $T=183120 221760 1 0 $X=182690 $Y=216640
X9113 1 2 199 226 BUJI3VX16 $T=332640 221760 0 180 $X=315970 $Y=216640
X9114 1 2 1014 180 BUJI3VX6 $T=37520 78400 1 180 $X=30370 $Y=77760
X9115 1 2 199 1269 BUJI3VX6 $T=309680 221760 1 0 $X=309250 $Y=216640
X9116 1 2 1009 87 86 1364 1435 ON31JI3VX1 $T=35840 69440 0 180 $X=30930 $Y=64320
X9117 1 2 90 270 274 251 1436 ON31JI3VX1 $T=47040 42560 0 180 $X=42130 $Y=37440
X9118 1 2 260 1022 261 1335 1298 ON31JI3VX1 $T=52080 203840 1 180 $X=47170 $Y=203200
X9119 1 2 343 342 347 1062 1437 ON31JI3VX1 $T=90160 212800 0 180 $X=85250 $Y=207680
X9120 1 2 426 873 136 418 1084 ON31JI3VX1 $T=144480 203840 1 180 $X=139570 $Y=203200
X9121 1 2 882 1231 136 874 1088 ON31JI3VX1 $T=152880 212800 0 180 $X=147970 $Y=207680
X9122 1 2 482 139 136 1096 1345 ON31JI3VX1 $T=166320 203840 1 180 $X=161410 $Y=203200
X9123 1 2 915 548 167 1349 1119 ON31JI3VX1 $T=223440 203840 1 180 $X=218530 $Y=203200
X9124 1 2 572 176 1122 592 1371 ON31JI3VX1 $T=231840 194880 0 0 $X=231410 $Y=194240
X9125 1 2 209 956 713 714 1324 ON31JI3VX1 $T=329280 203840 1 180 $X=324370 $Y=203200
X9126 1 2 734 713 1168 1278 1000 ON31JI3VX1 $T=332640 203840 0 0 $X=332210 $Y=203200
X9127 1 2 758 972 713 1203 1283 ON31JI3VX1 $T=344400 203840 1 0 $X=343970 $Y=198720
X9128 1 2 596 583 DLY4JI3VX1 $T=232960 212800 0 0 $X=232530 $Y=212160
X9129 1 2 SPI_CS 622 DLY4JI3VX1 $T=258720 221760 1 0 $X=258290 $Y=216640
X9130 1 2 131 151 180 NO2I1JI3VX2 $T=192640 42560 0 180 $X=187170 $Y=37440
X9131 1 2 199 643 BUJI3VX12 $T=275520 150080 1 0 $X=275090 $Y=144960
X9132 1 2 199 672 BUJI3VX12 $T=287840 150080 1 0 $X=287410 $Y=144960
X9133 1 2 648 up_switches<22> INJI3VX3 $T=281680 24640 1 0 $X=281250 $Y=19520
X9134 1 2 687 461 INJI3VX3 $T=304080 42560 1 0 $X=303650 $Y=37440
X9135 1 2 771 up_switches<3> INJI3VX3 $T=367360 24640 1 0 $X=366930 $Y=19520
X9136 1 2 776 up_switches<2> INJI3VX3 $T=370720 24640 1 0 $X=370290 $Y=19520
X9137 1 2 1438 1421 802 1021 987 NA4JI3VX0 $T=50400 60480 1 180 $X=46050 $Y=59840
X9138 1 2 858 1339 501 859 1439 NA4JI3VX0 $T=100800 185920 0 0 $X=100370 $Y=185280
X9139 1 2 1423 1197 1424 1135 1133 NA4JI3VX0 $T=255360 24640 0 0 $X=254930 $Y=24000
X9140 1 2 648 1198 776 771 664 NA4JI3VX0 $T=288960 24640 0 0 $X=288530 $Y=24000
X9141 1 2 959 518 1164 1360 1425 NA4JI3VX0 $T=329280 176960 1 180 $X=324930 $Y=176320
X9142 1 2 1215 1301 1393 355 OR3JI3VX1 $T=63840 194880 1 0 $X=63410 $Y=189760
X9143 1 2 630 934 682 1144 OR3JI3VX1 $T=272720 24640 1 0 $X=272290 $Y=19520
X9144 1 2 978 1178 1286 709 OR3JI3VX1 $T=349440 24640 1 180 $X=345090 $Y=24000
X9145 1 2 1144 664 1434 1197 NO3JI3VX1 $T=274960 24640 0 0 $X=274530 $Y=24000
X9146 1 2 1003 1333 240 436 277 FAJI3VX1 $T=23520 132160 0 0 $X=23090 $Y=131520
X9147 1 2 1002 1008 85 404 1333 FAJI3VX1 $T=23520 150080 0 0 $X=23090 $Y=149440
X9148 1 2 1005 1365 265 391 253 FAJI3VX1 $T=25200 105280 0 0 $X=24770 $Y=104640
X9149 1 2 790 1051 243 1016 1365 FAJI3VX1 $T=25200 114240 1 0 $X=24770 $Y=109120
X9150 1 2 809 1017 258 404 800 FAJI3VX1 $T=53760 150080 1 180 $X=38770 $Y=149440
X9151 1 2 1214 800 259 436 280 FAJI3VX1 $T=54320 150080 0 180 $X=39330 $Y=144960
X9152 1 2 95 805 100 391 1207 FAJI3VX1 $T=40880 114240 1 0 $X=40450 $Y=109120
X9153 1 2 97 290 812 1016 805 FAJI3VX1 $T=40880 114240 0 0 $X=40450 $Y=113600
X9154 1 2 294 272 265 1440 1026 FAJI3VX1 $T=41440 96320 0 0 $X=41010 $Y=95680
X9155 1 2 1366 1336 243 266 272 FAJI3VX1 $T=65520 105280 0 180 $X=50530 $Y=100160
X9156 1 2 1031 277 825 430 301 FAJI3VX1 $T=56560 132160 0 0 $X=56130 $Y=131520
X9157 1 2 103 315 823 393 290 FAJI3VX1 $T=58240 114240 0 0 $X=57810 $Y=113600
X9158 1 2 1032 280 298 430 101 FAJI3VX1 $T=58240 150080 1 0 $X=57810 $Y=144960
X9159 1 2 310 836 317 393 1051 FAJI3VX1 $T=68320 105280 0 0 $X=67890 $Y=104640
X9160 1 2 828 301 324 872 1055 FAJI3VX1 $T=70560 132160 1 0 $X=70130 $Y=127040
X9161 1 2 829 101 110 872 1056 FAJI3VX1 $T=70560 141120 1 0 $X=70130 $Y=136000
X9162 1 2 831 1056 106 1067 315 FAJI3VX1 $T=72800 123200 1 0 $X=72370 $Y=118080
X9163 1 2 1052 1055 331 1067 836 FAJI3VX1 $T=74480 114240 0 0 $X=74050 $Y=113600
X9164 1 2 921 188 BUJI3VX4 $T=233520 114240 0 180 $X=227490 $Y=109120
X9165 1 2 1306 489 INJI3VX1 $T=170800 185920 1 0 $X=170370 $Y=180800
X9166 1 2 553 549 INJI3VX1 $T=223440 221760 0 180 $X=221330 $Y=216640
X9167 1 2 549 246 DLY2JI3VX1 $T=175840 221760 1 0 $X=175410 $Y=216640
X9168 1 2 607 196 DLY2JI3VX1 $T=256480 212800 0 0 $X=256050 $Y=212160
X9169 1 2 269 256 246 104 84 269 SDFRRQJI3VX1 $T=42560 176960 1 180 $X=21970 $Y=176320
X9170 1 2 796 98 241 1015 94 98 SDFRRQJI3VX1 $T=43120 42560 1 180 $X=22530 $Y=41920
X9171 1 2 122 107 241 119 382 107 SDFRRQJI3VX1 $T=101360 60480 0 180 $X=80770 $Y=55360
X9172 1 2 122 350 241 402 382 350 SDFRRQJI3VX1 $T=101360 60480 1 180 $X=80770 $Y=59840
X9173 1 2 368 119 241 312 382 312 SDFRRQJI3VX1 $T=101360 69440 0 180 $X=80770 $Y=64320
X9174 1 2 368 118 241 348 382 348 SDFRRQJI3VX1 $T=101360 69440 1 180 $X=80770 $Y=68800
X9175 1 2 368 402 241 349 382 349 SDFRRQJI3VX1 $T=101360 78400 0 180 $X=80770 $Y=73280
X9176 1 2 121 356 241 402 382 356 SDFRRQJI3VX1 $T=105280 51520 1 180 $X=84690 $Y=50880
X9177 1 2 123 358 241 119 382 358 SDFRRQJI3VX1 $T=105280 132160 0 180 $X=84690 $Y=127040
X9178 1 2 123 359 241 402 382 359 SDFRRQJI3VX1 $T=105280 132160 1 180 $X=84690 $Y=131520
X9179 1 2 123 360 241 118 382 360 SDFRRQJI3VX1 $T=105280 141120 0 180 $X=84690 $Y=136000
X9180 1 2 123 109 241 364 382 109 SDFRRQJI3VX1 $T=105280 141120 1 180 $X=84690 $Y=140480
X9181 1 2 121 399 129 119 382 399 SDFRRQJI3VX1 $T=113120 60480 1 0 $X=112690 $Y=55360
X9182 1 2 121 400 129 118 382 400 SDFRRQJI3VX1 $T=113120 60480 0 0 $X=112690 $Y=59840
X9183 1 2 122 367 129 118 382 367 SDFRRQJI3VX1 $T=113120 69440 1 0 $X=112690 $Y=64320
X9184 1 2 122 411 132 396 382 411 SDFRRQJI3VX1 $T=113120 69440 0 0 $X=112690 $Y=68800
X9185 1 2 122 401 129 364 382 401 SDFRRQJI3VX1 $T=113120 87360 1 0 $X=112690 $Y=82240
X9186 1 2 382 118 129 402 188 118 SDFRRQJI3VX1 $T=113120 114240 0 0 $X=112690 $Y=113600
X9187 1 2 382 119 129 118 188 119 SDFRRQJI3VX1 $T=113120 123200 0 0 $X=112690 $Y=122560
X9188 1 2 382 402 129 364 188 402 SDFRRQJI3VX1 $T=113120 132160 1 0 $X=112690 $Y=127040
X9189 1 2 382 364 129 396 188 364 SDFRRQJI3VX1 $T=113120 132160 0 0 $X=112690 $Y=131520
X9190 1 2 382 396 129 454 188 396 SDFRRQJI3VX1 $T=113120 141120 1 0 $X=112690 $Y=136000
X9191 1 2 368 364 129 398 382 398 SDFRRQJI3VX1 $T=113120 141120 0 0 $X=112690 $Y=140480
X9192 1 2 123 403 129 454 382 403 SDFRRQJI3VX1 $T=113120 150080 1 0 $X=112690 $Y=144960
X9193 1 2 123 365 129 396 382 365 SDFRRQJI3VX1 $T=113120 159040 1 0 $X=112690 $Y=153920
X9194 1 2 368 396 129 408 382 408 SDFRRQJI3VX1 $T=115920 159040 0 0 $X=115490 $Y=158400
X9195 1 2 121 417 129 364 382 417 SDFRRQJI3VX1 $T=120960 78400 0 0 $X=120530 $Y=77760
X9196 1 2 121 432 132 396 382 432 SDFRRQJI3VX1 $T=125440 78400 1 0 $X=125010 $Y=73280
X9197 1 2 123 421 132 141 382 421 SDFRRQJI3VX1 $T=145600 96320 1 180 $X=125010 $Y=95680
X9198 1 2 368 454 129 397 382 397 SDFRRQJI3VX1 $T=125440 150080 0 0 $X=125010 $Y=149440
X9199 1 2 123 435 129 450 382 435 SDFRRQJI3VX1 $T=148400 96320 0 180 $X=127810 $Y=91200
X9200 1 2 368 141 132 447 382 447 SDFRRQJI3VX1 $T=153440 141120 1 180 $X=132850 $Y=140480
X9201 1 2 368 450 132 448 382 448 SDFRRQJI3VX1 $T=153440 150080 0 180 $X=132850 $Y=144960
X9202 1 2 382 450 129 141 188 450 SDFRRQJI3VX1 $T=133840 123200 0 0 $X=133410 $Y=122560
X9203 1 2 382 454 132 450 188 454 SDFRRQJI3VX1 $T=156240 132160 0 180 $X=135650 $Y=127040
X9204 1 2 121 471 132 450 382 471 SDFRRQJI3VX1 $T=142800 69440 0 0 $X=142370 $Y=68800
X9205 1 2 122 472 132 454 382 472 SDFRRQJI3VX1 $T=142800 87360 1 0 $X=142370 $Y=82240
X9206 1 2 121 475 132 454 382 475 SDFRRQJI3VX1 $T=145040 87360 0 0 $X=144610 $Y=86720
X9207 1 2 122 453 132 450 382 453 SDFRRQJI3VX1 $T=147280 78400 1 0 $X=146850 $Y=73280
X9208 1 2 123 427 132 488 382 427 SDFRRQJI3VX1 $T=167440 105280 0 180 $X=146850 $Y=100160
X9209 1 2 123 437 132 148 382 437 SDFRRQJI3VX1 $T=168560 96320 1 180 $X=147970 $Y=95680
X9210 1 2 368 148 132 458 382 458 SDFRRQJI3VX1 $T=175840 141120 1 180 $X=155250 $Y=140480
X9211 1 2 123 1090 132 138 382 1090 SDFRRQJI3VX1 $T=179200 114240 0 180 $X=158610 $Y=109120
X9212 1 2 382 146 147 138 188 146 SDFRRQJI3VX1 $T=159040 132160 1 0 $X=158610 $Y=127040
X9213 1 2 123 463 132 146 382 463 SDFRRQJI3VX1 $T=180320 105280 1 180 $X=159730 $Y=104640
X9214 1 2 382 488 147 146 188 488 SDFRRQJI3VX1 $T=160160 114240 0 0 $X=159730 $Y=113600
X9215 1 2 382 550 147 119 188 550 SDFRRQJI3VX1 $T=160160 123200 0 0 $X=159730 $Y=122560
X9216 1 2 196 148 132 488 188 148 SDFRRQJI3VX1 $T=180880 132160 1 180 $X=160290 $Y=131520
X9217 1 2 382 141 132 148 188 141 SDFRRQJI3VX1 $T=181440 141120 0 180 $X=160850 $Y=136000
X9218 1 2 368 488 132 492 SPI_CS 492 SDFRRQJI3VX1 $T=182000 150080 0 180 $X=161410 $Y=144960
X9219 1 2 368 146 147 503 SPI_CS 503 SDFRRQJI3VX1 $T=164080 150080 0 0 $X=163650 $Y=149440
X9220 1 2 121 508 147 141 SPI_CS 508 SDFRRQJI3VX1 $T=165200 78400 0 0 $X=164770 $Y=77760
X9221 1 2 122 509 147 141 SPI_CS 509 SDFRRQJI3VX1 $T=165760 87360 0 0 $X=165330 $Y=86720
X9222 1 2 122 510 147 148 SPI_CS 510 SDFRRQJI3VX1 $T=165760 96320 1 0 $X=165330 $Y=91200
X9223 1 2 121 143 147 148 SPI_CS 143 SDFRRQJI3VX1 $T=169680 123200 1 0 $X=169250 $Y=118080
X9224 1 2 368 138 147 495 SPI_CS 495 SDFRRQJI3VX1 $T=169680 159040 1 0 $X=169250 $Y=153920
X9225 1 2 121 517 147 488 SPI_CS 517 SDFRRQJI3VX1 $T=171360 96320 0 0 $X=170930 $Y=95680
X9226 1 2 122 1192 147 488 SPI_CS 1192 SDFRRQJI3VX1 $T=171360 105280 1 0 $X=170930 $Y=100160
X9227 1 2 121 1193 147 146 SPI_CS 1193 SDFRRQJI3VX1 $T=185920 87360 0 0 $X=185490 $Y=86720
X9228 1 2 123 512 147 547 SPI_CS 512 SDFRRQJI3VX1 $T=207200 150080 1 180 $X=186610 $Y=149440
X9229 1 2 122 533 147 146 SPI_CS 533 SDFRRQJI3VX1 $T=187600 96320 1 0 $X=187170 $Y=91200
X9230 1 2 121 157 147 550 SPI_CS 157 SDFRRQJI3VX1 $T=208320 105280 1 180 $X=187730 $Y=104640
X9231 1 2 122 160 147 550 SPI_CS 160 SDFRRQJI3VX1 $T=210000 123200 0 180 $X=189410 $Y=118080
X9232 1 2 368 197 147 149 SPI_CS 149 SDFRRQJI3VX1 $T=210000 159040 0 180 $X=189410 $Y=153920
X9233 1 2 123 535 147 550 SPI_CS 535 SDFRRQJI3VX1 $T=211120 132160 0 180 $X=190530 $Y=127040
X9234 1 2 121 168 568 577 SPI_CS 168 SDFRRQJI3VX1 $T=218960 87360 0 0 $X=218530 $Y=86720
X9235 1 2 122 574 568 577 SPI_CS 574 SDFRRQJI3VX1 $T=218960 96320 1 0 $X=218530 $Y=91200
X9236 1 2 121 575 568 547 SPI_CS 575 SDFRRQJI3VX1 $T=218960 96320 0 0 $X=218530 $Y=95680
X9237 1 2 122 169 568 547 SPI_CS 169 SDFRRQJI3VX1 $T=218960 105280 0 0 $X=218530 $Y=104640
X9238 1 2 368 224 584 576 SPI_CS 576 SDFRRQJI3VX1 $T=218960 114240 0 0 $X=218530 $Y=113600
X9239 1 2 196 577 568 547 188 577 SDFRRQJI3VX1 $T=218960 123200 1 0 $X=218530 $Y=118080
X9240 1 2 196 547 568 550 188 547 SDFRRQJI3VX1 $T=218960 123200 0 0 $X=218530 $Y=122560
X9241 1 2 196 138 568 554 188 138 SDFRRQJI3VX1 $T=218960 132160 1 0 $X=218530 $Y=127040
X9242 1 2 196 1128 568 577 188 1128 SDFRRQJI3VX1 $T=218960 132160 0 0 $X=218530 $Y=131520
X9243 1 2 368 644 568 551 SPI_CS 551 SDFRRQJI3VX1 $T=218960 141120 0 0 $X=218530 $Y=140480
X9244 1 2 368 616 568 552 SPI_CS 552 SDFRRQJI3VX1 $T=218960 150080 1 0 $X=218530 $Y=144960
X9245 1 2 123 573 568 1128 SPI_CS 573 SDFRRQJI3VX1 $T=218960 150080 0 0 $X=218530 $Y=149440
X9246 1 2 123 161 568 577 SPI_CS 161 SDFRRQJI3VX1 $T=218960 159040 1 0 $X=218530 $Y=153920
X9247 1 2 368 554 568 578 SPI_CS 578 SDFRRQJI3VX1 $T=218960 159040 0 0 $X=218530 $Y=158400
X9248 1 2 368 647 568 586 SPI_CS 586 SDFRRQJI3VX1 $T=246960 141120 0 180 $X=226370 $Y=136000
X9249 1 2 622 197 181 583 188 197 SDFRRQJI3VX1 $T=227360 221760 1 0 $X=226930 $Y=216640
X9250 1 2 122 175 568 591 SPI_CS 175 SDFRRQJI3VX1 $T=252000 105280 0 180 $X=231410 $Y=100160
X9251 1 2 368 662 568 571 SPI_CS 571 SDFRRQJI3VX1 $T=233520 114240 1 0 $X=233090 $Y=109120
X9252 1 2 123 597 568 591 SPI_CS 597 SDFRRQJI3VX1 $T=253680 168000 0 180 $X=233090 $Y=162880
X9253 1 2 121 610 568 1128 SPI_CS 610 SDFRRQJI3VX1 $T=239120 87360 0 0 $X=238690 $Y=86720
X9254 1 2 122 611 568 1128 SPI_CS 611 SDFRRQJI3VX1 $T=239120 96320 1 0 $X=238690 $Y=91200
X9255 1 2 123 923 584 603 SPI_CS 923 SDFRRQJI3VX1 $T=259280 150080 0 180 $X=238690 $Y=144960
X9256 1 2 368 683 568 579 SPI_CS 579 SDFRRQJI3VX1 $T=259280 150080 1 180 $X=238690 $Y=149440
X9257 1 2 123 183 584 608 SPI_CS 183 SDFRRQJI3VX1 $T=259280 159040 0 180 $X=238690 $Y=153920
X9258 1 2 121 614 584 591 SPI_CS 614 SDFRRQJI3VX1 $T=240240 105280 0 0 $X=239810 $Y=104640
X9259 1 2 368 195 568 580 SPI_CS 580 SDFRRQJI3VX1 $T=260400 114240 1 180 $X=239810 $Y=113600
X9260 1 2 368 773 568 581 SPI_CS 581 SDFRRQJI3VX1 $T=260400 123200 0 180 $X=239810 $Y=118080
X9261 1 2 368 719 568 606 SPI_CS 606 SDFRRQJI3VX1 $T=260400 123200 1 180 $X=239810 $Y=122560
X9262 1 2 196 608 181 1128 188 608 SDFRRQJI3VX1 $T=240800 132160 1 0 $X=240370 $Y=127040
X9263 1 2 196 603 181 608 188 603 SDFRRQJI3VX1 $T=261520 132160 1 180 $X=240930 $Y=131520
X9264 1 2 196 591 181 603 188 591 SDFRRQJI3VX1 $T=241920 141120 0 0 $X=241490 $Y=140480
X9265 1 2 196 624 181 1132 188 624 SDFRRQJI3VX1 $T=248080 212800 1 0 $X=247650 $Y=207680
X9266 1 2 122 625 568 608 SPI_CS 625 SDFRRQJI3VX1 $T=248640 87360 1 0 $X=248210 $Y=82240
X9267 1 2 121 626 568 603 SPI_CS 626 SDFRRQJI3VX1 $T=249200 78400 1 0 $X=248770 $Y=73280
X9268 1 2 122 627 568 603 SPI_CS 627 SDFRRQJI3VX1 $T=249200 78400 0 0 $X=248770 $Y=77760
X9269 1 2 121 628 568 608 SPI_CS 628 SDFRRQJI3VX1 $T=249200 96320 0 0 $X=248770 $Y=95680
X9270 1 2 196 1132 181 621 188 1132 SDFRRQJI3VX1 $T=269920 203840 0 180 $X=249330 $Y=198720
X9271 1 2 368 768 568 632 SPI_CS 632 SDFRRQJI3VX1 $T=253680 114240 1 0 $X=253250 $Y=109120
X9272 1 2 235 619 181 633 188 619 SDFRRQJI3VX1 $T=274960 168000 0 180 $X=254370 $Y=162880
X9273 1 2 196 1320 181 639 188 621 SDFRRQJI3VX1 $T=275520 194880 1 180 $X=254930 $Y=194240
X9274 1 2 196 633 181 637 188 633 SDFRRQJI3VX1 $T=276080 159040 1 180 $X=255490 $Y=158400
X9275 1 2 196 930 199 190 188 639 SDFRRQJI3VX1 $T=255920 194880 1 0 $X=255490 $Y=189760
X9276 1 2 196 1252 199 619 188 1142 SDFRRQJI3VX1 $T=257600 168000 0 0 $X=257170 $Y=167360
X9277 1 2 235 1258 181 1142 188 190 SDFRRQJI3VX1 $T=277760 176960 0 180 $X=257170 $Y=171840
X9278 1 2 123 615 584 637 SPI_CS 615 SDFRRQJI3VX1 $T=279440 159040 0 180 $X=258850 $Y=153920
X9279 1 2 121 193 584 637 SPI_CS 193 SDFRRQJI3VX1 $T=284480 105280 1 180 $X=263890 $Y=104640
X9280 1 2 196 773 181 224 188 773 SDFRRQJI3VX1 $T=264320 123200 1 0 $X=263890 $Y=118080
X9281 1 2 196 195 181 768 188 195 SDFRRQJI3VX1 $T=264320 123200 0 0 $X=263890 $Y=122560
X9282 1 2 196 637 181 591 188 637 SDFRRQJI3VX1 $T=264320 141120 1 0 $X=263890 $Y=136000
X9283 1 2 196 719 181 647 188 719 SDFRRQJI3VX1 $T=264880 132160 1 0 $X=264450 $Y=127040
X9284 1 2 235 647 181 616 188 647 SDFRRQJI3VX1 $T=264880 132160 0 0 $X=264450 $Y=131520
X9285 1 2 235 616 181 644 188 616 SDFRRQJI3VX1 $T=285600 141120 1 180 $X=265010 $Y=140480
X9286 1 2 122 654 584 138 235 654 SDFRRQJI3VX1 $T=269920 96320 0 0 $X=269490 $Y=95680
X9287 1 2 121 658 584 138 235 658 SDFRRQJI3VX1 $T=270480 96320 1 0 $X=270050 $Y=91200
X9288 1 2 122 660 219 616 235 660 SDFRRQJI3VX1 $T=272160 87360 1 0 $X=271730 $Y=82240
X9289 1 2 121 661 219 616 235 661 SDFRRQJI3VX1 $T=272160 87360 0 0 $X=271730 $Y=86720
X9290 1 2 123 675 219 616 235 675 SDFRRQJI3VX1 $T=277760 159040 0 0 $X=277330 $Y=158400
X9291 1 2 123 677 219 197 235 677 SDFRRQJI3VX1 $T=279440 159040 1 0 $X=279010 $Y=153920
X9292 1 2 235 768 219 662 188 768 SDFRRQJI3VX1 $T=288400 123200 1 0 $X=287970 $Y=118080
X9293 1 2 235 662 219 773 188 662 SDFRRQJI3VX1 $T=288400 123200 0 0 $X=287970 $Y=122560
X9294 1 2 235 683 219 195 188 683 SDFRRQJI3VX1 $T=288400 132160 1 0 $X=287970 $Y=127040
X9295 1 2 121 689 219 647 235 689 SDFRRQJI3VX1 $T=288960 78400 1 0 $X=288530 $Y=73280
X9296 1 2 121 690 219 197 235 690 SDFRRQJI3VX1 $T=288960 105280 0 0 $X=288530 $Y=104640
X9297 1 2 122 691 219 197 235 691 SDFRRQJI3VX1 $T=288960 114240 1 0 $X=288530 $Y=109120
X9298 1 2 235 224 219 719 188 224 SDFRRQJI3VX1 $T=288960 132160 0 0 $X=288530 $Y=131520
X9299 1 2 235 644 219 197 188 644 SDFRRQJI3VX1 $T=288960 141120 1 0 $X=288530 $Y=136000
X9300 1 2 235 554 219 683 188 554 SDFRRQJI3VX1 $T=309120 141120 1 180 $X=288530 $Y=140480
X9301 1 2 122 694 219 647 235 694 SDFRRQJI3VX1 $T=289520 78400 0 0 $X=289090 $Y=77760
X9302 1 2 123 203 219 647 235 203 SDFRRQJI3VX1 $T=289520 150080 0 0 $X=289090 $Y=149440
X9303 1 2 122 704 584 637 SPI_CS 704 SDFRRQJI3VX1 $T=292320 114240 0 0 $X=291890 $Y=113600
X9304 1 2 122 740 219 554 235 740 SDFRRQJI3VX1 $T=324800 69440 0 0 $X=324370 $Y=68800
X9305 1 2 121 741 219 554 235 741 SDFRRQJI3VX1 $T=324800 78400 1 0 $X=324370 $Y=73280
X9306 1 2 121 742 219 683 235 742 SDFRRQJI3VX1 $T=324800 87360 1 0 $X=324370 $Y=82240
X9307 1 2 122 213 219 683 235 213 SDFRRQJI3VX1 $T=324800 87360 0 0 $X=324370 $Y=86720
X9308 1 2 121 716 219 644 235 716 SDFRRQJI3VX1 $T=324800 114240 0 0 $X=324370 $Y=113600
X9309 1 2 122 718 219 644 235 718 SDFRRQJI3VX1 $T=324800 123200 1 0 $X=324370 $Y=118080
X9310 1 2 121 739 199 719 235 739 SDFRRQJI3VX1 $T=324800 123200 0 0 $X=324370 $Y=122560
X9311 1 2 123 743 219 644 235 743 SDFRRQJI3VX1 $T=324800 132160 1 0 $X=324370 $Y=127040
X9312 1 2 123 214 219 683 235 214 SDFRRQJI3VX1 $T=324800 150080 1 0 $X=324370 $Y=144960
X9313 1 2 123 720 199 554 235 720 SDFRRQJI3VX1 $T=326480 159040 1 0 $X=326050 $Y=153920
X9314 1 2 122 751 199 224 235 751 SDFRRQJI3VX1 $T=336560 114240 1 0 $X=336130 $Y=109120
X9315 1 2 123 752 199 719 235 752 SDFRRQJI3VX1 $T=336560 132160 0 0 $X=336130 $Y=131520
X9316 1 2 123 748 199 224 235 748 SDFRRQJI3VX1 $T=336560 141120 1 0 $X=336130 $Y=136000
X9317 1 2 121 755 199 224 235 755 SDFRRQJI3VX1 $T=337120 105280 0 0 $X=336690 $Y=104640
X9318 1 2 121 759 219 195 235 759 SDFRRQJI3VX1 $T=338240 78400 0 0 $X=337810 $Y=77760
X9319 1 2 122 757 219 195 235 757 SDFRRQJI3VX1 $T=338240 96320 1 0 $X=337810 $Y=91200
X9320 1 2 121 770 199 773 235 770 SDFRRQJI3VX1 $T=344960 123200 1 0 $X=344530 $Y=118080
X9321 1 2 122 1182 199 719 235 1182 SDFRRQJI3VX1 $T=344960 123200 0 0 $X=344530 $Y=122560
X9322 1 2 123 231 199 195 235 231 SDFRRQJI3VX1 $T=344960 132160 1 0 $X=344530 $Y=127040
X9323 1 2 121 782 199 662 235 782 SDFRRQJI3VX1 $T=360640 96320 0 0 $X=360210 $Y=95680
X9324 1 2 122 783 199 662 235 783 SDFRRQJI3VX1 $T=360640 105280 1 0 $X=360210 $Y=100160
X9325 1 2 121 784 199 768 235 784 SDFRRQJI3VX1 $T=360640 114240 1 0 $X=360210 $Y=109120
X9326 1 2 122 233 199 768 235 233 SDFRRQJI3VX1 $T=360640 114240 0 0 $X=360210 $Y=113600
X9327 1 2 123 785 199 662 235 785 SDFRRQJI3VX1 $T=360640 132160 0 0 $X=360210 $Y=131520
X9328 1 2 123 786 199 768 235 786 SDFRRQJI3VX1 $T=360640 141120 1 0 $X=360210 $Y=136000
X9329 1 2 123 775 199 773 235 775 SDFRRQJI3VX1 $T=360640 141120 0 0 $X=360210 $Y=140480
X9330 1 2 122 232 199 773 235 232 SDFRRQJI3VX1 $T=365120 123200 1 0 $X=364690 $Y=118080
X9331 1 2 129 241 BUJI3VX3 $T=100800 168000 1 0 $X=100370 $Y=162880
X9332 1 2 1078 enable BUJI3VX3 $T=122640 185920 0 0 $X=122210 $Y=185280
X9333 1 2 151 687 BUJI3VX3 $T=192640 24640 0 0 $X=192210 $Y=24000
X9334 1 2 199 938 BUJI3VX3 $T=280000 168000 0 0 $X=279570 $Y=167360
X9335 1 2 199 650 BUJI3VX3 $T=280560 168000 1 0 $X=280130 $Y=162880
X9336 1 2 1095 up_switches<18> BUJI3VX3 $T=295680 24640 0 0 $X=295250 $Y=24000
X9337 1 2 199 1263 BUJI3VX3 $T=295680 176960 1 0 $X=295250 $Y=171840
X9338 1 2 671 up_switches<17> BUJI3VX3 $T=299040 24640 1 0 $X=298610 $Y=19520
X9339 1 2 199 943 BUJI3VX3 $T=301280 212800 1 0 $X=300850 $Y=207680
X9340 1 2 682 up_switches<16> BUJI3VX3 $T=302960 24640 1 0 $X=302530 $Y=19520
X9341 1 2 199 697 BUJI3VX3 $T=302960 212800 0 0 $X=302530 $Y=212160
X9342 1 2 199 949 BUJI3VX3 $T=303520 150080 1 0 $X=303090 $Y=144960
X9343 1 2 199 1160 BUJI3VX3 $T=306880 176960 1 0 $X=306450 $Y=171840
X9344 1 2 688 up_switches<15> BUJI3VX3 $T=307440 24640 1 0 $X=307010 $Y=19520
X9345 1 2 701 up_switches<14> BUJI3VX3 $T=311360 24640 1 0 $X=310930 $Y=19520
X9346 1 2 199 712 BUJI3VX3 $T=313600 203840 0 0 $X=313170 $Y=203200
X9347 1 2 532 up_switches<13> BUJI3VX3 $T=327600 24640 0 180 $X=323250 $Y=19520
X9348 1 2 715 up_switches<12> BUJI3VX3 $T=337120 24640 1 180 $X=332770 $Y=24000
X9349 1 2 199 733 BUJI3VX3 $T=334880 159040 0 0 $X=334450 $Y=158400
X9350 1 2 736 up_switches<11> BUJI3VX3 $T=341040 24640 0 180 $X=336690 $Y=19520
X9351 1 2 1166 up_switches<10> BUJI3VX3 $T=341040 24640 1 180 $X=336690 $Y=24000
X9352 1 2 976 up_switches<9> BUJI3VX3 $T=344960 24640 1 180 $X=340610 $Y=24000
X9353 1 2 977 up_switches<8> BUJI3VX3 $T=348880 24640 0 180 $X=344530 $Y=19520
X9354 1 2 1178 up_switches<7> BUJI3VX3 $T=352800 24640 0 180 $X=348450 $Y=19520
X9355 1 2 1286 up_switches<6> BUJI3VX3 $T=352240 24640 0 0 $X=351810 $Y=24000
X9356 1 2 750 up_switches<5> BUJI3VX3 $T=353360 24640 1 0 $X=352930 $Y=19520
X9357 1 2 199 1289 BUJI3VX3 $T=355040 203840 0 0 $X=354610 $Y=203200
X9358 1 2 199 983 BUJI3VX3 $T=358960 203840 0 0 $X=358530 $Y=203200
X9359 1 2 767 up_switches<4> BUJI3VX3 $T=364560 24640 1 180 $X=360210 $Y=24000
X9360 1 2 215 up_switches<1> BUJI3VX3 $T=374080 24640 1 0 $X=373650 $Y=19520
X9361 1 2 204 up_switches<0> BUJI3VX3 $T=379120 24640 1 0 $X=378690 $Y=19520
X9362 1 2 247 87 INJI3VX0 $T=29120 69440 1 0 $X=28690 $Y=64320
X9363 1 2 1013 1205 INJI3VX0 $T=39200 69440 1 0 $X=38770 $Y=64320
X9364 1 2 104 261 INJI3VX0 $T=44240 194880 1 180 $X=42130 $Y=194240
X9365 1 2 1022 797 INJI3VX0 $T=47040 203840 0 180 $X=44930 $Y=198720
X9366 1 2 1009 1422 INJI3VX0 $T=47600 60480 1 0 $X=47170 $Y=55360
X9367 1 2 93 801 INJI3VX0 $T=49840 42560 1 180 $X=47730 $Y=41920
X9368 1 2 90 804 INJI3VX0 $T=49840 42560 0 0 $X=49410 $Y=41920
X9369 1 2 1210 1438 INJI3VX0 $T=52640 60480 1 180 $X=50530 $Y=59840
X9370 1 2 1024 1028 INJI3VX0 $T=52080 185920 1 0 $X=51650 $Y=180800
X9371 1 2 89 292 INJI3VX0 $T=53200 194880 1 0 $X=52770 $Y=189760
X9372 1 2 305 270 INJI3VX0 $T=57680 33600 1 180 $X=55570 $Y=32960
X9373 1 2 278 263 INJI3VX0 $T=59360 51520 0 180 $X=57250 $Y=46400
X9374 1 2 276 1440 INJI3VX0 $T=59360 96320 1 180 $X=57250 $Y=95680
X9375 1 2 341 266 INJI3VX0 $T=59360 105280 1 180 $X=57250 $Y=104640
X9376 1 2 98 815 INJI3VX0 $T=58240 42560 1 0 $X=57810 $Y=37440
X9377 1 2 279 1414 INJI3VX0 $T=59920 185920 1 0 $X=59490 $Y=180800
X9378 1 2 297 1034 INJI3VX0 $T=63840 176960 1 180 $X=61730 $Y=176320
X9379 1 2 105 1441 INJI3VX0 $T=64400 203840 1 180 $X=62290 $Y=203200
X9380 1 2 1037 1043 INJI3VX0 $T=64400 212800 1 0 $X=63970 $Y=207680
X9381 1 2 293 826 INJI3VX0 $T=68320 203840 1 0 $X=67890 $Y=198720
X9382 1 2 308 1053 INJI3VX0 $T=75040 194880 1 0 $X=74610 $Y=189760
X9383 1 2 344 108 INJI3VX0 $T=81760 105280 0 180 $X=79650 $Y=100160
X9384 1 2 324 1070 INJI3VX0 $T=83440 123200 0 0 $X=83010 $Y=122560
X9385 1 2 335 322 INJI3VX0 $T=85680 194880 1 180 $X=83570 $Y=194240
X9386 1 2 336 835 INJI3VX0 $T=91280 203840 0 180 $X=89170 $Y=198720
X9387 1 2 113 112 INJI3VX0 $T=91840 96320 1 180 $X=89730 $Y=95680
X9388 1 2 342 1222 INJI3VX0 $T=92400 212800 1 0 $X=91970 $Y=207680
X9389 1 2 991 267 INJI3VX0 $T=95200 203840 1 180 $X=93090 $Y=203200
X9390 1 2 853 327 INJI3VX0 $T=96880 176960 1 180 $X=94770 $Y=176320
X9391 1 2 296 347 INJI3VX0 $T=95200 203840 0 0 $X=94770 $Y=203200
X9392 1 2 345 1075 INJI3VX0 $T=98000 105280 1 0 $X=97570 $Y=100160
X9393 1 2 1223 858 INJI3VX0 $T=100240 185920 1 0 $X=99810 $Y=180800
X9394 1 2 856 1397 INJI3VX0 $T=113120 24640 1 0 $X=112690 $Y=19520
X9395 1 2 379 1077 INJI3VX0 $T=124320 194880 0 180 $X=122210 $Y=189760
X9396 1 2 115 1079 INJI3VX0 $T=128800 33600 1 180 $X=126690 $Y=32960
X9397 1 2 863 414 INJI3VX0 $T=133840 194880 0 0 $X=133410 $Y=194240
X9398 1 2 413 868 INJI3VX0 $T=137760 24640 1 180 $X=135650 $Y=24000
X9399 1 2 426 1083 INJI3VX0 $T=137760 194880 1 180 $X=135650 $Y=194240
X9400 1 2 412 873 INJI3VX0 $T=137200 203840 0 0 $X=136770 $Y=203200
X9401 1 2 452 876 INJI3VX0 $T=142800 194880 0 0 $X=142370 $Y=194240
X9402 1 2 442 875 INJI3VX0 $T=149520 33600 1 180 $X=147410 $Y=32960
X9403 1 2 446 879 INJI3VX0 $T=148960 24640 0 0 $X=148530 $Y=24000
X9404 1 2 882 451 INJI3VX0 $T=151760 194880 0 0 $X=151330 $Y=194240
X9405 1 2 425 136 INJI3VX0 $T=155120 203840 1 180 $X=153010 $Y=203200
X9406 1 2 1305 1233 INJI3VX0 $T=155680 185920 1 0 $X=155250 $Y=180800
X9407 1 2 887 1092 INJI3VX0 $T=159600 24640 1 180 $X=157490 $Y=24000
X9408 1 2 886 1094 INJI3VX0 $T=157920 203840 1 0 $X=157490 $Y=198720
X9409 1 2 481 1101 INJI3VX0 $T=163520 24640 0 0 $X=163090 $Y=24000
X9410 1 2 482 477 INJI3VX0 $T=166320 194880 1 180 $X=164210 $Y=194240
X9411 1 2 496 1102 INJI3VX0 $T=171920 194880 1 180 $X=169810 $Y=194240
X9412 1 2 137 897 INJI3VX0 $T=175280 24640 0 0 $X=174850 $Y=24000
X9413 1 2 150 1104 INJI3VX0 $T=182000 194880 1 180 $X=179890 $Y=194240
X9414 1 2 900 1398 INJI3VX0 $T=184240 33600 0 180 $X=182130 $Y=28480
X9415 1 2 518 307 INJI3VX0 $T=184240 194880 0 180 $X=182130 $Y=189760
X9416 1 2 511 1399 INJI3VX0 $T=188160 24640 0 180 $X=186050 $Y=19520
X9417 1 2 1108 502 INJI3VX0 $T=188720 203840 0 180 $X=186610 $Y=198720
X9418 1 2 527 152 INJI3VX0 $T=190960 212800 0 0 $X=190530 $Y=212160
X9419 1 2 528 1239 INJI3VX0 $T=193760 212800 0 0 $X=193330 $Y=212160
X9420 1 2 903 1400 INJI3VX0 $T=198240 33600 1 180 $X=196130 $Y=32960
X9421 1 2 910 1401 INJI3VX0 $T=201040 24640 0 180 $X=198930 $Y=19520
X9422 1 2 167 159 INJI3VX0 $T=201040 203840 0 180 $X=198930 $Y=198720
X9423 1 2 541 912 INJI3VX0 $T=201040 203840 1 0 $X=200610 $Y=198720
X9424 1 2 1113 908 INJI3VX0 $T=204400 203840 0 180 $X=202290 $Y=198720
X9425 1 2 917 1310 INJI3VX0 $T=218960 42560 1 0 $X=218530 $Y=37440
X9426 1 2 174 914 INJI3VX0 $T=221200 24640 1 180 $X=219090 $Y=24000
X9427 1 2 560 1118 INJI3VX0 $T=221200 42560 1 0 $X=220770 $Y=37440
X9428 1 2 557 556 INJI3VX0 $T=227360 185920 1 180 $X=225250 $Y=185280
X9429 1 2 1126 1123 INJI3VX0 $T=233520 24640 1 180 $X=231410 $Y=24000
X9430 1 2 570 176 INJI3VX0 $T=236880 203840 1 180 $X=234770 $Y=203200
X9431 1 2 594 1372 INJI3VX0 $T=240240 194880 0 180 $X=238130 $Y=189760
X9432 1 2 572 925 INJI3VX0 $T=240240 194880 1 0 $X=239810 $Y=189760
X9433 1 2 588 1420 INJI3VX0 $T=246960 194880 1 0 $X=246530 $Y=189760
X9434 1 2 926 1402 INJI3VX0 $T=248640 33600 1 0 $X=248210 $Y=28480
X9435 1 2 927 929 INJI3VX0 $T=250880 42560 0 0 $X=250450 $Y=41920
X9436 1 2 194 1319 INJI3VX0 $T=266000 42560 1 0 $X=265570 $Y=37440
X9437 1 2 636 1257 INJI3VX0 $T=272160 33600 1 0 $X=271730 $Y=28480
X9438 1 2 enable 126 INJI3VX0 $T=276080 185920 0 0 $X=275650 $Y=185280
X9439 1 2 196 657 INJI3VX0 $T=277760 194880 1 0 $X=277330 $Y=189760
X9440 1 2 659 674 INJI3VX0 $T=281120 221760 1 0 $X=280690 $Y=216640
X9441 1 2 940 1403 INJI3VX0 $T=286160 33600 0 180 $X=284050 $Y=28480
X9442 1 2 1149 1262 INJI3VX0 $T=287280 42560 1 0 $X=286850 $Y=37440
X9443 1 2 1152 944 INJI3VX0 $T=299600 33600 0 0 $X=299170 $Y=32960
X9444 1 2 942 696 INJI3VX0 $T=301280 185920 0 0 $X=300850 $Y=185280
X9445 1 2 700 1153 INJI3VX0 $T=301280 194880 1 0 $X=300850 $Y=189760
X9446 1 2 1158 951 INJI3VX0 $T=306320 33600 1 0 $X=305890 $Y=28480
X9447 1 2 703 206 INJI3VX0 $T=313600 185920 1 0 $X=313170 $Y=180800
X9448 1 2 1411 202 INJI3VX0 $T=315840 203840 0 180 $X=313730 $Y=198720
X9449 1 2 708 713 INJI3VX0 $T=324800 194880 0 0 $X=324370 $Y=194240
X9450 1 2 1163 1404 INJI3VX0 $T=328160 42560 0 180 $X=326050 $Y=37440
X9451 1 2 734 722 INJI3VX0 $T=328160 194880 1 180 $X=326050 $Y=194240
X9452 1 2 222 957 INJI3VX0 $T=328720 51520 1 0 $X=328290 $Y=46400
X9453 1 2 721 958 INJI3VX0 $T=330960 203840 1 0 $X=330530 $Y=198720
X9454 1 2 1168 1361 INJI3VX0 $T=334320 203840 0 180 $X=332210 $Y=198720
X9455 1 2 1171 1405 INJI3VX0 $T=335440 33600 0 180 $X=333330 $Y=28480
X9456 1 2 220 1280 INJI3VX0 $T=337680 185920 1 0 $X=337250 $Y=180800
X9457 1 2 965 1172 INJI3VX0 $T=337680 194880 1 0 $X=337250 $Y=189760
X9458 1 2 1279 1173 INJI3VX0 $T=338800 42560 1 0 $X=338370 $Y=37440
X9459 1 2 971 735 INJI3VX0 $T=341040 168000 1 180 $X=338930 $Y=167360
X9460 1 2 968 1406 INJI3VX0 $T=341040 24640 1 0 $X=340610 $Y=19520
X9461 1 2 975 973 INJI3VX0 $T=346640 168000 1 180 $X=344530 $Y=167360
X9462 1 2 761 979 INJI3VX0 $T=350560 42560 1 0 $X=350130 $Y=37440
X9463 1 2 1179 738 INJI3VX0 $T=355040 194880 0 180 $X=352930 $Y=189760
X9464 1 2 981 1330 INJI3VX0 $T=356720 176960 0 0 $X=356290 $Y=176320
X9465 1 2 758 1001 INJI3VX0 $T=357840 185920 0 0 $X=357410 $Y=185280
X9466 1 2 1290 1183 INJI3VX0 $T=364560 24640 0 0 $X=364130 $Y=24000
X9467 1 2 228 1407 INJI3VX0 $T=370720 33600 0 180 $X=368610 $Y=28480
X9468 1 2 1009 1435 1013 NA2JI3VX0 $T=36960 69440 1 0 $X=36530 $Y=64320
X9469 1 2 252 1011 794 NA2JI3VX0 $T=42000 60480 1 180 $X=39330 $Y=59840
X9470 1 2 1385 1010 795 NA2JI3VX0 $T=43680 203840 0 180 $X=41010 $Y=198720
X9471 1 2 263 1021 252 NA2JI3VX0 $T=47040 60480 0 180 $X=44370 $Y=55360
X9472 1 2 254 1436 1186 NA2JI3VX0 $T=49840 42560 0 180 $X=47170 $Y=37440
X9473 1 2 1209 1298 795 NA2JI3VX0 $T=50400 203840 0 180 $X=47730 $Y=198720
X9474 1 2 89 1022 1025 NA2JI3VX0 $T=53200 194880 1 180 $X=50530 $Y=194240
X9475 1 2 283 802 87 NA2JI3VX0 $T=56560 69440 0 180 $X=53890 $Y=64320
X9476 1 2 96 271 1422 NA2JI3VX0 $T=58800 60480 0 180 $X=56130 $Y=55360
X9477 1 2 322 1299 260 NA2JI3VX0 $T=59360 203840 0 180 $X=56690 $Y=198720
X9478 1 2 1040 814 334 NA2JI3VX0 $T=63840 87360 1 180 $X=61170 $Y=86720
X9479 1 2 1217 818 334 NA2JI3VX0 $T=67760 87360 1 180 $X=65090 $Y=86720
X9480 1 2 823 1218 327 NA2JI3VX0 $T=68880 105280 0 180 $X=66210 $Y=100160
X9481 1 2 314 822 334 NA2JI3VX0 $T=71120 87360 1 180 $X=68450 $Y=86720
X9482 1 2 293 833 308 NA2JI3VX0 $T=71120 203840 0 0 $X=70690 $Y=203200
X9483 1 2 1045 300 292 NA2JI3VX0 $T=73920 194880 0 180 $X=71250 $Y=189760
X9484 1 2 1219 832 334 NA2JI3VX0 $T=75600 87360 1 180 $X=72930 $Y=86720
X9485 1 2 303 1057 1053 NA2JI3VX0 $T=73360 185920 1 0 $X=72930 $Y=180800
X9486 1 2 337 1442 334 NA2JI3VX0 $T=77840 96320 1 0 $X=77410 $Y=91200
X9487 1 2 106 1302 327 NA2JI3VX0 $T=85120 114240 1 0 $X=84690 $Y=109120
X9488 1 2 110 845 327 NA2JI3VX0 $T=89600 123200 1 180 $X=86930 $Y=122560
X9489 1 2 343 1437 1068 NA2JI3VX0 $T=90160 212800 1 0 $X=89730 $Y=207680
X9490 1 2 1221 1443 334 NA2JI3VX0 $T=92960 96320 0 180 $X=90290 $Y=91200
X9491 1 2 127 1439 854 NA2JI3VX0 $T=99680 185920 1 180 $X=97010 $Y=185280
X9492 1 2 330 1337 1068 NA2JI3VX0 $T=98560 203840 0 0 $X=98130 $Y=203200
X9493 1 2 856 1374 180 NA2JI3VX0 $T=99680 24640 1 0 $X=99250 $Y=19520
X9494 1 2 1188 1076 131 NA2JI3VX0 $T=102480 24640 0 0 $X=102050 $Y=24000
X9495 1 2 enable 859 336 NA2JI3VX0 $T=102480 203840 0 0 $X=102050 $Y=203200
X9496 1 2 1188 1224 180 NA2JI3VX0 $T=113680 24640 0 0 $X=113250 $Y=24000
X9497 1 2 379 124 1368 NA2JI3VX0 $T=118160 194880 0 180 $X=115490 $Y=189760
X9498 1 2 1077 372 1368 NA2JI3VX0 $T=121520 194880 0 180 $X=118850 $Y=189760
X9499 1 2 376 1227 180 NA2JI3VX0 $T=123200 24640 0 0 $X=122770 $Y=24000
X9500 1 2 379 514 1226 NA2JI3VX0 $T=123200 203840 1 0 $X=122770 $Y=198720
X9501 1 2 376 1426 131 NA2JI3VX0 $T=127120 24640 0 0 $X=126690 $Y=24000
X9502 1 2 115 1228 180 NA2JI3VX0 $T=128800 33600 1 0 $X=128370 $Y=28480
X9503 1 2 865 867 180 NA2JI3VX0 $T=133280 24640 0 0 $X=132850 $Y=24000
X9504 1 2 407 1082 1444 NA2JI3VX0 $T=134960 203840 1 0 $X=134530 $Y=198720
X9505 1 2 865 1427 131 NA2JI3VX0 $T=135520 33600 1 0 $X=135090 $Y=28480
X9506 1 2 1085 434 414 NA2JI3VX0 $T=136640 185920 1 0 $X=136210 $Y=180800
X9507 1 2 413 871 180 NA2JI3VX0 $T=138320 24640 0 0 $X=137890 $Y=24000
X9508 1 2 409 440 1083 NA2JI3VX0 $T=138320 185920 0 0 $X=137890 $Y=185280
X9509 1 2 869 1084 1444 NA2JI3VX0 $T=138320 203840 1 0 $X=137890 $Y=198720
X9510 1 2 1086 992 180 NA2JI3VX0 $T=139440 33600 0 0 $X=139010 $Y=32960
X9511 1 2 431 1229 180 NA2JI3VX0 $T=141680 24640 0 0 $X=141250 $Y=24000
X9512 1 2 1086 1428 131 NA2JI3VX0 $T=143360 33600 0 0 $X=142930 $Y=32960
X9513 1 2 434 1304 1419 NA2JI3VX0 $T=146160 185920 1 0 $X=145730 $Y=180800
X9514 1 2 442 457 180 NA2JI3VX0 $T=150640 33600 0 0 $X=150210 $Y=32960
X9515 1 2 467 1232 180 NA2JI3VX0 $T=154000 24640 0 0 $X=153570 $Y=24000
X9516 1 2 884 1305 451 NA2JI3VX0 $T=156240 194880 0 180 $X=153570 $Y=189760
X9517 1 2 886 1231 135 NA2JI3VX0 $T=154000 194880 0 0 $X=153570 $Y=194240
X9518 1 2 1097 1235 180 NA2JI3VX0 $T=162960 33600 1 0 $X=162530 $Y=28480
X9519 1 2 476 888 477 NA2JI3VX0 $T=164640 185920 1 0 $X=164210 $Y=180800
X9520 1 2 1099 485 180 NA2JI3VX0 $T=165200 24640 0 0 $X=164770 $Y=24000
X9521 1 2 1102 891 425 NA2JI3VX0 $T=170240 194880 1 180 $X=167570 $Y=194240
X9522 1 2 515 470 1102 NA2JI3VX0 $T=168560 185920 1 0 $X=168130 $Y=180800
X9523 1 2 899 1105 180 NA2JI3VX0 $T=179200 33600 0 0 $X=178770 $Y=32960
X9524 1 2 507 1107 180 NA2JI3VX0 $T=185360 24640 1 180 $X=182690 $Y=24000
X9525 1 2 528 538 527 NA2JI3VX0 $T=187040 212800 0 0 $X=186610 $Y=212160
X9526 1 2 904 1369 180 NA2JI3VX0 $T=197120 42560 0 180 $X=194450 $Y=37440
X9527 1 2 1309 1112 180 NA2JI3VX0 $T=198800 24640 1 180 $X=196130 $Y=24000
X9528 1 2 904 1114 131 NA2JI3VX0 $T=201040 42560 1 0 $X=200610 $Y=37440
X9529 1 2 903 909 180 NA2JI3VX0 $T=201600 33600 0 0 $X=201170 $Y=32960
X9530 1 2 559 531 908 NA2JI3VX0 $T=205520 194880 1 0 $X=205090 $Y=189760
X9531 1 2 561 1313 180 NA2JI3VX0 $T=210560 24640 1 180 $X=207890 $Y=24000
X9532 1 2 1120 1115 180 NA2JI3VX0 $T=210560 33600 1 180 $X=207890 $Y=32960
X9533 1 2 174 1315 180 NA2JI3VX0 $T=221760 33600 1 0 $X=221330 $Y=28480
X9534 1 2 915 1119 558 NA2JI3VX0 $T=225680 203840 1 180 $X=223010 $Y=203200
X9535 1 2 561 1430 542 NA2JI3VX0 $T=225120 24640 0 0 $X=224690 $Y=24000
X9536 1 2 1120 918 542 NA2JI3VX0 $T=225680 33600 0 0 $X=225250 $Y=32960
X9537 1 2 557 1352 915 NA2JI3VX0 $T=227920 203840 1 180 $X=225250 $Y=203200
X9538 1 2 917 1243 180 NA2JI3VX0 $T=226240 42560 1 0 $X=225810 $Y=37440
X9539 1 2 919 1117 180 NA2JI3VX0 $T=232400 42560 0 180 $X=229730 $Y=37440
X9540 1 2 1125 1242 180 NA2JI3VX0 $T=232960 24640 0 180 $X=230290 $Y=19520
X9541 1 2 560 1247 180 NA2JI3VX0 $T=232400 33600 0 0 $X=231970 $Y=32960
X9542 1 2 582 1371 1248 NA2JI3VX0 $T=233520 203840 1 0 $X=233090 $Y=198720
X9543 1 2 919 1127 542 NA2JI3VX0 $T=236320 42560 0 180 $X=233650 $Y=37440
X9544 1 2 1125 1431 542 NA2JI3VX0 $T=234640 24640 1 0 $X=234210 $Y=19520
X9545 1 2 172 170 556 NA2JI3VX0 $T=238560 194880 0 180 $X=235890 $Y=189760
X9546 1 2 1126 1354 180 NA2JI3VX0 $T=238560 24640 0 0 $X=238130 $Y=24000
X9547 1 2 589 1433 542 NA2JI3VX0 $T=240240 42560 1 0 $X=239810 $Y=37440
X9548 1 2 589 1249 180 NA2JI3VX0 $T=241360 33600 0 0 $X=240930 $Y=32960
X9549 1 2 1410 602 1432 NA2JI3VX0 $T=245840 203840 1 0 $X=245410 $Y=198720
X9550 1 2 926 1355 180 NA2JI3VX0 $T=248080 42560 1 0 $X=247650 $Y=37440
X9551 1 2 598 594 1420 NA2JI3VX0 $T=252000 194880 0 180 $X=249330 $Y=189760
X9552 1 2 928 1131 180 NA2JI3VX0 $T=252000 42560 1 0 $X=251570 $Y=37440
X9553 1 2 927 1317 180 NA2JI3VX0 $T=254240 42560 0 0 $X=253810 $Y=41920
X9554 1 2 928 1318 542 NA2JI3VX0 $T=258160 42560 0 180 $X=255490 $Y=37440
X9555 1 2 623 1136 542 NA2JI3VX0 $T=262640 42560 0 180 $X=259970 $Y=37440
X9556 1 2 194 1138 180 NA2JI3VX0 $T=263760 33600 1 180 $X=261090 $Y=32960
X9557 1 2 623 1255 180 NA2JI3VX0 $T=263760 33600 0 0 $X=263330 $Y=32960
X9558 1 2 633 1137 192 NA2JI3VX0 $T=263760 150080 0 0 $X=263330 $Y=149440
X9559 1 2 932 1139 198 NA2JI3VX0 $T=269360 33600 0 0 $X=268930 $Y=32960
X9560 1 2 1146 1145 1143 NA2JI3VX0 $T=280000 203840 0 180 $X=277330 $Y=198720
X9561 1 2 1260 1321 198 NA2JI3VX0 $T=278880 33600 0 0 $X=278450 $Y=32960
X9562 1 2 668 1261 198 NA2JI3VX0 $T=295120 33600 1 180 $X=292450 $Y=32960
X9563 1 2 676 1264 198 NA2JI3VX0 $T=299040 33600 1 180 $X=296370 $Y=32960
X9564 1 2 1155 692 1153 NA2JI3VX0 $T=300720 185920 1 0 $X=300290 $Y=180800
X9565 1 2 945 1267 198 NA2JI3VX0 $T=304080 33600 0 0 $X=303650 $Y=32960
X9566 1 2 700 956 705 NA2JI3VX0 $T=310800 185920 1 0 $X=310370 $Y=180800
X9567 1 2 727 1378 198 NA2JI3VX0 $T=316400 33600 1 180 $X=313730 $Y=32960
X9568 1 2 725 212 198 NA2JI3VX0 $T=325360 51520 1 0 $X=324930 $Y=46400
X9569 1 2 961 717 958 NA2JI3VX0 $T=325360 185920 0 0 $X=324930 $Y=185280
X9570 1 2 209 1324 998 NA2JI3VX0 $T=327600 203840 0 180 $X=324930 $Y=198720
X9571 1 2 721 1273 1274 NA2JI3VX0 $T=328160 194880 0 0 $X=327730 $Y=194240
X9572 1 2 717 960 1165 NA2JI3VX0 $T=329280 185920 1 0 $X=328850 $Y=180800
X9573 1 2 962 999 198 NA2JI3VX0 $T=330400 33600 0 0 $X=329970 $Y=32960
X9574 1 2 223 1379 198 NA2JI3VX0 $T=333760 33600 0 180 $X=331090 $Y=28480
X9575 1 2 225 1326 198 NA2JI3VX0 $T=335440 42560 1 0 $X=335010 $Y=37440
X9576 1 2 734 1000 1274 NA2JI3VX0 $T=337680 203840 0 180 $X=335010 $Y=198720
X9577 1 2 744 220 1172 NA2JI3VX0 $T=341040 185920 1 180 $X=338370 $Y=185280
X9578 1 2 974 971 973 NA2JI3VX0 $T=344400 168000 1 180 $X=341730 $Y=167360
X9579 1 2 981 972 1176 NA2JI3VX0 $T=346640 185920 1 180 $X=343970 $Y=185280
X9580 1 2 758 1283 1281 NA2JI3VX0 $T=346080 194880 0 0 $X=345650 $Y=194240
X9581 1 2 229 1284 198 NA2JI3VX0 $T=350000 42560 0 180 $X=347330 $Y=37440
X9582 1 2 230 730 760 NA2JI3VX0 $T=351120 176960 0 180 $X=348450 $Y=171840
X9583 1 2 982 766 198 NA2JI3VX0 $T=357840 24640 0 0 $X=357410 $Y=24000
X9584 1 2 1412 1291 198 NA2JI3VX0 $T=359520 33600 0 0 $X=359090 $Y=32960
X9585 1 2 1181 230 1001 NA2JI3VX0 $T=365120 176960 0 180 $X=362450 $Y=171840
X9586 1 2 104 1005 256 265 1296 AO22JI3VX1 $T=31360 105280 0 180 $X=25890 $Y=100160
X9587 1 2 1003 104 256 240 237 AO22JI3VX1 $T=28560 132160 1 0 $X=28130 $Y=127040
X9588 1 2 1002 104 256 85 238 AO22JI3VX1 $T=29120 150080 1 0 $X=28690 $Y=144960
X9589 1 2 791 104 256 1334 239 AO22JI3VX1 $T=29120 168000 0 0 $X=28690 $Y=167360
X9590 1 2 104 790 256 243 793 AO22JI3VX1 $T=29680 114240 0 0 $X=29250 $Y=113600
X9591 1 2 104 244 256 88 242 AO22JI3VX1 $T=33040 105280 1 0 $X=32610 $Y=100160
X9592 1 2 1445 104 256 289 250 AO22JI3VX1 $T=45360 185920 1 180 $X=39890 $Y=185280
X9593 1 2 1446 104 256 89 792 AO22JI3VX1 $T=45360 194880 0 180 $X=39890 $Y=189760
X9594 1 2 1208 104 256 279 249 AO22JI3VX1 $T=47040 176960 0 180 $X=41570 $Y=171840
X9595 1 2 809 296 267 258 248 AO22JI3VX1 $T=49280 159040 0 180 $X=43810 $Y=153920
X9596 1 2 1214 296 267 259 799 AO22JI3VX1 $T=49840 141120 1 180 $X=44370 $Y=140480
X9597 1 2 1297 296 267 803 806 AO22JI3VX1 $T=45920 168000 1 0 $X=45490 $Y=162880
X9598 1 2 296 1185 267 91 1018 AO22JI3VX1 $T=52640 123200 1 180 $X=47170 $Y=122560
X9599 1 2 296 95 267 100 1019 AO22JI3VX1 $T=55440 123200 0 180 $X=49970 $Y=118080
X9600 1 2 1037 1441 296 1418 268 AO22JI3VX1 $T=61600 203840 1 180 $X=56130 $Y=203200
X9601 1 2 1032 296 267 298 817 AO22JI3VX1 $T=57680 150080 0 0 $X=57250 $Y=149440
X9602 1 2 296 97 267 812 1216 AO22JI3VX1 $T=58240 123200 1 0 $X=57810 $Y=118080
X9603 1 2 296 103 267 823 287 AO22JI3VX1 $T=70560 123200 0 180 $X=65090 $Y=118080
X9604 1 2 1031 104 256 825 304 AO22JI3VX1 $T=69440 141120 0 0 $X=69010 $Y=140480
X9605 1 2 104 310 256 317 299 AO22JI3VX1 $T=78960 114240 0 180 $X=73490 $Y=109120
X9606 1 2 831 296 267 106 352 AO22JI3VX1 $T=73920 123200 0 0 $X=73490 $Y=122560
X9607 1 2 829 296 267 110 346 AO22JI3VX1 $T=74480 150080 1 0 $X=74050 $Y=144960
X9608 1 2 828 104 256 324 316 AO22JI3VX1 $T=76160 141120 0 0 $X=75730 $Y=140480
X9609 1 2 1058 296 267 326 329 AO22JI3VX1 $T=76160 203840 0 0 $X=75730 $Y=203200
X9610 1 2 505 313 835 enable 256 AO22JI3VX1 $T=83440 194880 1 180 $X=77970 $Y=194240
X9611 1 2 1052 104 256 331 351 AO22JI3VX1 $T=79520 114240 1 0 $X=79090 $Y=109120
X9612 1 2 392 425 420 863 380 AO22JI3VX1 $T=128240 203840 1 180 $X=122770 $Y=203200
X9613 1 2 505 1080 374 enable 420 AO22JI3VX1 $T=123760 194880 0 0 $X=123330 $Y=194240
X9614 1 2 467 151 180 887 1095 AO22JI3VX1 $T=156240 33600 1 0 $X=155810 $Y=28480
X9615 1 2 1097 151 180 481 671 AO22JI3VX1 $T=167440 33600 1 0 $X=167010 $Y=28480
X9616 1 2 1099 151 180 137 682 AO22JI3VX1 $T=170240 24640 0 0 $X=169810 $Y=24000
X9617 1 2 899 151 180 900 688 AO22JI3VX1 $T=180880 42560 1 0 $X=180450 $Y=37440
X9618 1 2 507 151 180 511 701 AO22JI3VX1 $T=187600 24640 0 0 $X=187170 $Y=24000
X9619 1 2 1309 687 180 910 532 AO22JI3VX1 $T=201600 24640 0 0 $X=201170 $Y=24000
X9620 1 2 537 159 912 528 529 AO22JI3VX1 $T=208880 203840 1 180 $X=203410 $Y=203200
X9621 1 2 1116 159 912 1113 913 AO22JI3VX1 $T=204960 203840 1 0 $X=204530 $Y=198720
X9622 1 2 557 558 159 1350 916 AO22JI3VX1 $T=225120 203840 0 180 $X=219650 $Y=198720
X9623 1 2 932 687 198 636 715 AO22JI3VX1 $T=272160 33600 0 0 $X=271730 $Y=32960
X9624 1 2 676 687 198 1152 204 AO22JI3VX1 $T=297920 42560 1 0 $X=297490 $Y=37440
X9625 1 2 945 687 198 1158 736 AO22JI3VX1 $T=308000 33600 0 0 $X=307570 $Y=32960
X9626 1 2 955 708 998 703 210 AO22JI3VX1 $T=316960 194880 0 180 $X=311490 $Y=189760
X9627 1 2 727 687 198 1163 215 AO22JI3VX1 $T=324800 33600 0 0 $X=324370 $Y=32960
X9628 1 2 725 687 198 222 1166 AO22JI3VX1 $T=325920 42560 0 0 $X=325490 $Y=41920
X9629 1 2 962 687 198 1171 767 AO22JI3VX1 $T=335440 33600 1 0 $X=335010 $Y=28480
X9630 1 2 708 964 965 126 746 AO22JI3VX1 $T=336000 194880 0 0 $X=335570 $Y=194240
X9631 1 2 223 687 198 968 750 AO22JI3VX1 $T=341600 33600 1 0 $X=341170 $Y=28480
X9632 1 2 225 687 198 1279 976 AO22JI3VX1 $T=341600 42560 1 0 $X=341170 $Y=37440
X9633 1 2 708 1373 1281 1285 1202 AO22JI3VX1 $T=348880 194880 0 0 $X=348450 $Y=194240
X9634 1 2 1447 708 975 126 774 AO22JI3VX1 $T=350560 176960 0 0 $X=350130 $Y=176320
X9635 1 2 1177 708 981 126 1292 AO22JI3VX1 $T=350560 185920 0 0 $X=350130 $Y=185280
X9636 1 2 1412 687 198 228 1178 AO22JI3VX1 $T=357840 33600 1 180 $X=352370 $Y=32960
X9637 1 2 982 687 198 1290 1286 AO22JI3VX1 $T=358400 33600 0 180 $X=352930 $Y=28480
X9638 1 2 229 687 198 761 977 AO22JI3VX1 $T=358400 42560 0 180 $X=352930 $Y=37440
X9639 1 2 709 1271 706 698 1198 OR4JI3VX2 $T=316960 24640 1 180 $X=309250 $Y=24000
X9640 1 2 489 132 INJI3VX2 $T=173600 168000 1 0 $X=173170 $Y=162880
X9641 1 2 489 147 INJI3VX2 $T=177520 185920 0 0 $X=177090 $Y=185280
X9642 1 2 185 640 INJI3VX2 $T=223440 221760 1 0 $X=223010 $Y=216640
X9643 1 2 180 798 257 1204 AO21JI3VX1 $T=43120 78400 1 180 $X=38210 $Y=77760
X9644 1 2 104 1022 256 795 AO21JI3VX1 $T=49840 194880 1 180 $X=44930 $Y=194240
X9645 1 2 308 267 830 1041 AO21JI3VX1 $T=73360 212800 0 180 $X=68450 $Y=207680
X9646 1 2 848 1070 345 1303 AO21JI3VX1 $T=92400 114240 0 180 $X=87490 $Y=109120
X9647 1 2 873 425 420 1444 AO21JI3VX1 $T=145040 203840 0 180 $X=140130 $Y=198720
X9648 1 2 126 680 1151 1150 AO21JI3VX1 $T=296800 194880 0 180 $X=291890 $Y=189760
X9649 1 2 288 1039 339 NO2I1JI3VX1 $T=64960 194880 0 0 $X=64530 $Y=194240
X9650 1 2 1057 311 1415 NO2I1JI3VX1 $T=77840 176960 1 180 $X=74050 $Y=176320
X9651 1 2 383 1049 317 NO2I1JI3VX1 $T=80080 96320 1 180 $X=76290 $Y=95680
X9652 1 2 111 357 331 NO2I1JI3VX1 $T=86800 105280 0 0 $X=86370 $Y=104640
X9653 1 2 333 847 343 NO2I1JI3VX1 $T=88480 185920 0 0 $X=88050 $Y=185280
X9654 1 2 339 851 1071 NO2I1JI3VX1 $T=91840 194880 0 0 $X=91410 $Y=194240
X9655 1 2 1226 336 379 NO2I1JI3VX1 $T=122080 203840 0 180 $X=118290 $Y=198720
X9656 1 2 369 1226 116 NO2I1JI3VX1 $T=123200 194880 1 180 $X=119410 $Y=194240
X9657 1 2 407 130 864 NO2I1JI3VX1 $T=128800 185920 0 0 $X=128370 $Y=185280
X9658 1 2 405 410 130 NO2I1JI3VX1 $T=134400 194880 1 0 $X=133970 $Y=189760
X9659 1 2 891 898 420 NO2I1JI3VX1 $T=166880 203840 1 0 $X=166450 $Y=198720
X9660 1 2 153 1417 528 NO2I1JI3VX1 $T=196560 194880 0 0 $X=196130 $Y=194240
X9661 1 2 171 536 915 NO2I1JI3VX1 $T=222320 185920 1 180 $X=218530 $Y=185280
X9662 1 2 192 1141 633 NO2I1JI3VX1 $T=267120 150080 0 0 $X=266690 $Y=149440
X9663 1 2 692 947 1159 NO2I1JI3VX1 $T=306320 176960 1 180 $X=302530 $Y=176320
X9664 1 2 296 989 826 308 NA3JI3VX0 $T=70000 194880 0 0 $X=69570 $Y=194240
X9665 1 2 832 1044 1396 1218 NA3JI3VX0 $T=74480 96320 1 180 $X=71250 $Y=95680
X9666 1 2 320 838 837 333 NA3JI3VX0 $T=81200 185920 1 0 $X=80770 $Y=180800
X9667 1 2 1442 1060 839 1302 NA3JI3VX0 $T=83440 96320 1 0 $X=83010 $Y=91200
X9668 1 2 340 114 338 333 NA3JI3VX0 $T=85680 185920 1 0 $X=85250 $Y=180800
X9669 1 2 1443 1066 846 845 NA3JI3VX0 $T=89600 96320 0 180 $X=86370 $Y=91200
X9670 1 2 1077 374 369 116 NA3JI3VX0 $T=115920 194880 0 0 $X=115490 $Y=194240
X9671 1 2 480 462 440 1189 NA3JI3VX0 $T=149520 194880 0 180 $X=146290 $Y=189760
X9672 1 2 1091 373 1448 1089 NA3JI3VX0 $T=155120 185920 1 180 $X=151890 $Y=185280
X9673 1 2 410 1376 470 474 NA3JI3VX0 $T=160160 194880 1 0 $X=159730 $Y=189760
X9674 1 2 889 466 1448 888 NA3JI3VX0 $T=164080 185920 1 180 $X=160850 $Y=185280
X9675 1 2 1449 1191 888 890 NA3JI3VX0 $T=167440 185920 1 180 $X=164210 $Y=185280
X9676 1 2 1429 889 890 474 NA3JI3VX0 $T=167440 194880 0 180 $X=164210 $Y=189760
X9677 1 2 425 1236 502 496 NA3JI3VX0 $T=172480 194880 0 0 $X=172050 $Y=194240
X9678 1 2 1108 139 496 150 NA3JI3VX0 $T=179200 194880 1 180 $X=175970 $Y=194240
X9679 1 2 1377 221 953 200 NA3JI3VX0 $T=310800 176960 1 0 $X=310370 $Y=171840
X9680 1 2 708 1268 202 680 NA3JI3VX0 $T=313600 194880 1 180 $X=310370 $Y=194240
X9681 1 2 711 954 731 953 NA3JI3VX0 $T=316960 176960 0 180 $X=313730 $Y=171840
X9682 1 2 221 1325 1162 731 NA3JI3VX0 $T=333200 176960 0 0 $X=332770 $Y=176320
X9683 1 2 180 257 1012 OR2JI3VX0 $T=43120 69440 1 180 $X=39330 $Y=68800
X9684 1 2 252 263 987 OR2JI3VX0 $T=41440 60480 1 0 $X=41010 $Y=55360
X9685 1 2 1043 824 1050 OR2JI3VX0 $T=69440 185920 0 0 $X=69010 $Y=185280
X9686 1 2 833 1043 1061 OR2JI3VX0 $T=74480 203840 1 0 $X=74050 $Y=198720
X9687 1 2 1083 409 1189 OR2JI3VX0 $T=138320 194880 1 0 $X=137890 $Y=189760
X9688 1 2 477 476 890 OR2JI3VX0 $T=161280 185920 1 0 $X=160850 $Y=180800
X9689 1 2 1104 493 474 OR2JI3VX0 $T=180880 194880 0 180 $X=177090 $Y=189760
X9690 1 2 514 126 501 OR2JI3VX0 $T=184800 185920 1 180 $X=181010 $Y=185280
X9691 1 2 1239 902 906 OR2JI3VX0 $T=193200 194880 0 0 $X=192770 $Y=194240
X9692 1 2 176 1129 1353 OR2JI3VX0 $T=235760 185920 0 180 $X=231970 $Y=180800
X9693 1 2 1153 1155 200 OR2JI3VX0 $T=296800 176960 0 0 $X=296370 $Y=176320
X9694 1 2 970 738 967 OR2JI3VX0 $T=343280 194880 0 180 $X=339490 $Y=189760
X9695 1 2 enable 1341 127 321 1225 AO211JI3VX1 $T=113120 185920 0 0 $X=112690 $Y=185280
X9696 1 2 791 295 245 1008 HAJI3VX1 $T=28000 159040 0 0 $X=27570 $Y=158400
X9697 1 2 1297 295 262 1017 HAJI3VX1 $T=48160 159040 1 180 $X=39890 $Y=158400
X9698 1 2 1208 269 279 1024 HAJI3VX1 $T=44800 176960 0 0 $X=44370 $Y=176320
X9699 1 2 1445 289 1024 1025 HAJI3VX1 $T=45920 185920 0 0 $X=45490 $Y=185280
X9700 1 2 392 863 866 412 HAJI3VX1 $T=126000 203840 1 0 $X=125570 $Y=198720
X9701 1 2 1147 663 1450 1143 HAJI3VX1 $T=281120 203840 1 0 $X=280690 $Y=198720
X9702 1 2 673 669 1322 1450 HAJI3VX1 $T=296800 203840 0 180 $X=288530 $Y=198720
X9703 1 2 1447 975 1175 1176 HAJI3VX1 $T=349440 176960 1 180 $X=341170 $Y=176320
X9704 1 2 843 850 851 353 OA21JI3VX1 $T=91280 194880 1 0 $X=90850 $Y=189760
X9705 1 2 1145 1143 936 1140 OA21JI3VX1 $T=276640 203840 0 180 $X=271730 $Y=198720
X9706 1 2 89 1025 1446 EO2JI3VX0 $T=52080 194880 0 180 $X=46050 $Y=189760
X9707 1 2 1054 344 1065 EO2JI3VX0 $T=81760 105280 1 0 $X=81330 $Y=100160
X9708 1 2 345 855 990 EO2JI3VX0 $T=96880 105280 0 180 $X=90850 $Y=100160
X9709 1 2 624 IC_addr<1> 1134 EO2JI3VX0 $T=250880 212800 0 0 $X=250450 $Y=212160
X9710 1 2 1132 IC_addr<0> 931 EO2JI3VX0 $T=253120 221760 1 0 $X=252690 $Y=216640
X9711 1 2 981 1176 1177 EO2JI3VX0 $T=345520 185920 1 0 $X=345090 $Y=180800
X9712 1 2 838 854 842 1220 NO3JI3VX0 $T=84560 185920 0 0 $X=84130 $Y=185280
X9713 1 2 1416 334 1223 321 NO3JI3VX0 $T=101360 176960 1 180 $X=97570 $Y=176320
X9714 1 2 444 1089 1419 881 NO3JI3VX0 $T=148400 185920 1 0 $X=147970 $Y=180800
X9715 1 2 462 1091 1376 1191 NO3JI3VX0 $T=156800 194880 1 0 $X=156370 $Y=189760
X9716 1 2 1238 1111 536 153 NO3JI3VX0 $T=196000 185920 1 180 $X=192210 $Y=185280
X9717 1 2 1134 192 931 634 NO3JI3VX0 $T=259840 203840 0 0 $X=259410 $Y=203200
X9718 1 2 1165 1360 1170 724 NO3JI3VX0 $T=330960 185920 1 180 $X=327170 $Y=185280
X9719 1 2 969 966 227 126 NO3JI3VX0 $T=342160 176960 0 180 $X=338370 $Y=171840
X9720 1 2 847 338 340 849 335 AN31JI3VX1 $T=90720 185920 1 0 $X=90290 $Y=180800
X9721 1 2 1384 1111 565 321 501 AN31JI3VX1 $T=189840 185920 1 180 $X=185490 $Y=185280
X9722 1 2 1413 1021 798 AND2JI3VX0 $T=48160 69440 0 180 $X=44370 $Y=64320
X9723 1 2 445 452 866 AND2JI3VX0 $T=142800 194880 1 180 $X=139010 $Y=194240
X9724 1 2 152 902 153 AND2JI3VX0 $T=193200 194880 0 180 $X=189410 $Y=189760
X9725 1 2 176 1129 566 AND2JI3VX0 $T=239120 185920 0 180 $X=235330 $Y=180800
X9726 1 2 659 656 1322 AND2JI3VX0 $T=291760 212800 0 180 $X=287970 $Y=207680
X9727 1 2 1246 565 922 1394 NO3I1JI3VX1 $T=236880 185920 1 180 $X=231970 $Y=185280
X9728 1 2 1093 1094 1448 1233 460 AN211JI3VX1 $T=160160 185920 1 180 $X=155250 $Y=185280
X9729 1 2 1276 206 1162 735 749 AN211JI3VX1 $T=335440 168000 1 180 $X=330530 $Y=167360
X9730 1 2 745 738 1164 1280 218 AN211JI3VX1 $T=340480 176960 1 180 $X=335570 $Y=176320
X9731 1 2 1102 515 1449 896 NO22JI3VX1 $T=168560 185920 0 0 $X=168130 $Y=185280
X9732 1 2 619 121 1141 NA2JI3VX2 $T=275520 150080 0 180 $X=271170 $Y=144960
X9733 1 2 619 1137 368 NO2JI3VX2 $T=259280 150080 0 0 $X=258850 $Y=149440
X9734 1 2 1137 122 619 NA2I1JI3VX2 $T=262080 150080 1 0 $X=261650 $Y=144960
X9735 1 2 619 123 1141 NA2I1JI3VX2 $T=273280 150080 0 0 $X=272850 $Y=149440
X9736 1 2 DECAP25JI3V $T=20160 24640 1 0 $X=19730 $Y=19520
X9737 1 2 DECAP25JI3V $T=20160 24640 0 0 $X=19730 $Y=24000
X9738 1 2 DECAP25JI3V $T=20160 87360 0 0 $X=19730 $Y=86720
X9739 1 2 DECAP25JI3V $T=20160 168000 1 0 $X=19730 $Y=162880
X9740 1 2 DECAP25JI3V $T=20160 212800 0 0 $X=19730 $Y=212160
X9741 1 2 DECAP25JI3V $T=20160 221760 1 0 $X=19730 $Y=216640
X9742 1 2 DECAP25JI3V $T=33040 33600 1 0 $X=32610 $Y=28480
X9743 1 2 DECAP25JI3V $T=34160 24640 1 0 $X=33730 $Y=19520
X9744 1 2 DECAP25JI3V $T=34160 87360 0 0 $X=33730 $Y=86720
X9745 1 2 DECAP25JI3V $T=34160 221760 1 0 $X=33730 $Y=216640
X9746 1 2 DECAP25JI3V $T=47040 33600 1 0 $X=46610 $Y=28480
X9747 1 2 DECAP25JI3V $T=99120 123200 0 0 $X=98690 $Y=122560
X9748 1 2 DECAP25JI3V $T=191520 96320 0 0 $X=191090 $Y=95680
X9749 1 2 DECAP25JI3V $T=212240 105280 1 0 $X=211810 $Y=100160
X9750 1 2 DECAP25JI3V $T=213920 114240 1 0 $X=213490 $Y=109120
X9751 1 2 DECAP25JI3V $T=260400 114240 0 0 $X=259970 $Y=113600
X9752 1 2 DECAP25JI3V $T=301280 69440 0 0 $X=300850 $Y=68800
X9753 1 2 DECAP25JI3V $T=309120 132160 0 0 $X=308690 $Y=131520
X9754 1 2 DECAP25JI3V $T=310800 78400 0 0 $X=310370 $Y=77760
X9755 1 2 DECAP25JI3V $T=341040 221760 1 0 $X=340610 $Y=216640
X9756 1 2 DECAP25JI3V $T=344400 212800 0 0 $X=343970 $Y=212160
X9757 1 2 DECAP25JI3V $T=344960 87360 1 0 $X=344530 $Y=82240
X9758 1 2 DECAP25JI3V $T=344960 212800 1 0 $X=344530 $Y=207680
X9759 1 2 DECAP25JI3V $T=355040 221760 1 0 $X=354610 $Y=216640
X9760 1 2 DECAP25JI3V $T=358400 105280 0 0 $X=357970 $Y=104640
X9761 1 2 DECAP25JI3V $T=358400 212800 0 0 $X=357970 $Y=212160
X9762 1 2 DECAP25JI3V $T=358960 87360 1 0 $X=358530 $Y=82240
X9763 1 2 DECAP25JI3V $T=358960 212800 1 0 $X=358530 $Y=207680
X9764 1 2 DECAP25JI3V $T=361760 150080 1 0 $X=361330 $Y=144960
X9765 1 2 DECAP25JI3V $T=362880 203840 0 0 $X=362450 $Y=203200
X9766 1 2 DECAP25JI3V $T=364000 176960 0 0 $X=363570 $Y=176320
X9767 1 2 DECAP25JI3V $T=365120 132160 1 0 $X=364690 $Y=127040
X9768 1 2 DECAP25JI3V $T=366240 24640 0 0 $X=365810 $Y=24000
X9769 1 2 DECAP25JI3V $T=367360 203840 1 0 $X=366930 $Y=198720
X9770 1 2 DECAP25JI3V $T=369040 221760 1 0 $X=368610 $Y=216640
X9771 1 2 DECAP25JI3V $T=371280 194880 0 0 $X=370850 $Y=194240
X9772 1 2 DECAP25JI3V $T=372400 105280 0 0 $X=371970 $Y=104640
X9773 1 2 DECAP25JI3V $T=372400 194880 1 0 $X=371970 $Y=189760
X9774 1 2 DECAP25JI3V $T=372400 212800 0 0 $X=371970 $Y=212160
X9775 1 2 DECAP25JI3V $T=372960 87360 1 0 $X=372530 $Y=82240
X9776 1 2 DECAP25JI3V $T=372960 212800 1 0 $X=372530 $Y=207680
X9777 1 2 DECAP25JI3V $T=374080 185920 1 0 $X=373650 $Y=180800
X9778 1 2 DECAP25JI3V $T=374640 185920 0 0 $X=374210 $Y=185280
X9779 1 2 DECAP25JI3V $T=375200 123200 0 0 $X=374770 $Y=122560
X9780 1 2 DECAP25JI3V $T=375760 150080 1 0 $X=375330 $Y=144960
X9781 1 2 DECAP25JI3V $T=376880 203840 0 0 $X=376450 $Y=203200
X9782 1 2 DECAP25JI3V $T=378000 176960 0 0 $X=377570 $Y=176320
X9783 1 2 DECAP25JI3V $T=378560 78400 0 0 $X=378130 $Y=77760
X9784 1 2 DECAP25JI3V $T=392560 87360 1 180 $X=378130 $Y=86720
X9785 1 2 DECAP25JI3V $T=378560 96320 1 0 $X=378130 $Y=91200
X9786 1 2 DECAP25JI3V $T=378560 150080 0 0 $X=378130 $Y=149440
X9787 1 2 DECAP25JI3V $T=379120 51520 1 0 $X=378690 $Y=46400
X9788 1 2 DECAP25JI3V $T=379120 51520 0 0 $X=378690 $Y=50880
X9789 1 2 DECAP25JI3V $T=379120 60480 1 0 $X=378690 $Y=55360
X9790 1 2 DECAP25JI3V $T=379120 60480 0 0 $X=378690 $Y=59840
X9791 1 2 DECAP25JI3V $T=379120 69440 0 0 $X=378690 $Y=68800
X9792 1 2 DECAP25JI3V $T=379120 132160 1 0 $X=378690 $Y=127040
X9793 1 2 DECAP25JI3V $T=379120 159040 0 0 $X=378690 $Y=158400
X9794 1 2 DECAP25JI3V $T=379120 168000 0 0 $X=378690 $Y=167360
X9795 1 2 DECAP25JI3V $T=379680 33600 0 0 $X=379250 $Y=32960
X9796 1 2 DECAP25JI3V $T=380240 24640 0 0 $X=379810 $Y=24000
X9797 1 2 DECAP25JI3V $T=380240 159040 1 0 $X=379810 $Y=153920
X9798 1 2 DECAP25JI3V $T=380800 33600 1 0 $X=380370 $Y=28480
X9799 1 2 DECAP25JI3V $T=380800 114240 1 0 $X=380370 $Y=109120
X9800 1 2 DECAP25JI3V $T=380800 141120 0 0 $X=380370 $Y=140480
X9801 1 2 DECAP25JI3V $T=381360 203840 1 0 $X=380930 $Y=198720
X9802 1 2 DECAP25JI3V $T=381920 96320 0 0 $X=381490 $Y=95680
X9803 1 2 DECAP25JI3V $T=381920 105280 1 0 $X=381490 $Y=100160
X9804 1 2 DECAP25JI3V $T=381920 114240 0 0 $X=381490 $Y=113600
X9805 1 2 DECAP25JI3V $T=381920 132160 0 0 $X=381490 $Y=131520
X9806 1 2 DECAP25JI3V $T=381920 141120 1 0 $X=381490 $Y=136000
X9807 1 2 DECAP25JI3V $T=382480 69440 1 0 $X=382050 $Y=64320
X9808 1 2 DECAP25JI3V $T=383040 24640 1 0 $X=382610 $Y=19520
X9809 1 2 DECAP25JI3V $T=383040 221760 1 0 $X=382610 $Y=216640
X9810 1 2 DECAP25JI3V $T=385280 194880 0 0 $X=384850 $Y=194240
X9811 1 2 DECAP25JI3V $T=386400 105280 0 0 $X=385970 $Y=104640
X9812 1 2 DECAP25JI3V $T=386400 123200 1 0 $X=385970 $Y=118080
X9813 1 2 DECAP25JI3V $T=386400 194880 1 0 $X=385970 $Y=189760
X9814 1 2 DECAP25JI3V $T=386400 212800 0 0 $X=385970 $Y=212160
X9815 1 2 DECAP25JI3V $T=386960 78400 1 0 $X=386530 $Y=73280
X9816 1 2 DECAP25JI3V $T=386960 87360 1 0 $X=386530 $Y=82240
X9817 1 2 DECAP25JI3V $T=386960 212800 1 0 $X=386530 $Y=207680
X9818 1 2 DECAP25JI3V $T=387520 176960 1 0 $X=387090 $Y=171840
X9819 1 2 DECAP25JI3V $T=388080 185920 1 0 $X=387650 $Y=180800
X9820 1 2 DECAP25JI3V $T=388640 185920 0 0 $X=388210 $Y=185280
X9821 1 2 DECAP25JI3V $T=389200 123200 0 0 $X=388770 $Y=122560
X9822 1 2 DECAP25JI3V $T=389760 150080 1 0 $X=389330 $Y=144960
X9823 1 2 DECAP25JI3V $T=390880 203840 0 0 $X=390450 $Y=203200
X9824 1 2 DECAP25JI3V $T=392000 176960 0 0 $X=391570 $Y=176320
X9825 1 2 DECAP25JI3V $T=392560 78400 0 0 $X=392130 $Y=77760
X9826 1 2 DECAP25JI3V $T=392560 87360 0 0 $X=392130 $Y=86720
X9827 1 2 DECAP25JI3V $T=392560 96320 1 0 $X=392130 $Y=91200
X9828 1 2 DECAP25JI3V $T=392560 150080 0 0 $X=392130 $Y=149440
X9829 1 2 DECAP25JI3V $T=393120 42560 1 0 $X=392690 $Y=37440
X9830 1 2 DECAP25JI3V $T=393120 42560 0 0 $X=392690 $Y=41920
X9831 1 2 DECAP25JI3V $T=393120 51520 1 0 $X=392690 $Y=46400
X9832 1 2 DECAP25JI3V $T=393120 51520 0 0 $X=392690 $Y=50880
X9833 1 2 DECAP25JI3V $T=393120 60480 1 0 $X=392690 $Y=55360
X9834 1 2 DECAP25JI3V $T=393120 60480 0 0 $X=392690 $Y=59840
X9835 1 2 DECAP25JI3V $T=393120 69440 0 0 $X=392690 $Y=68800
X9836 1 2 DECAP25JI3V $T=393120 132160 1 0 $X=392690 $Y=127040
X9837 1 2 DECAP25JI3V $T=393120 159040 0 0 $X=392690 $Y=158400
X9838 1 2 DECAP25JI3V $T=393120 168000 1 0 $X=392690 $Y=162880
X9839 1 2 DECAP25JI3V $T=393120 168000 0 0 $X=392690 $Y=167360
X9840 1 2 DECAP25JI3V $T=393680 33600 0 0 $X=393250 $Y=32960
X9841 1 2 DECAP25JI3V $T=394240 24640 0 0 $X=393810 $Y=24000
X9842 1 2 DECAP25JI3V $T=394240 159040 1 0 $X=393810 $Y=153920
X9843 1 2 DECAP25JI3V $T=394800 33600 1 0 $X=394370 $Y=28480
X9844 1 2 DECAP25JI3V $T=394800 114240 1 0 $X=394370 $Y=109120
X9845 1 2 DECAP25JI3V $T=394800 141120 0 0 $X=394370 $Y=140480
X9846 1 2 DECAP25JI3V $T=395360 203840 1 0 $X=394930 $Y=198720
X9847 1 2 DECAP25JI3V $T=395920 96320 0 0 $X=395490 $Y=95680
X9848 1 2 DECAP25JI3V $T=395920 105280 1 0 $X=395490 $Y=100160
X9849 1 2 DECAP25JI3V $T=395920 114240 0 0 $X=395490 $Y=113600
X9850 1 2 DECAP25JI3V $T=395920 132160 0 0 $X=395490 $Y=131520
X9851 1 2 DECAP25JI3V $T=395920 141120 1 0 $X=395490 $Y=136000
X9852 1 2 DECAP25JI3V $T=396480 69440 1 0 $X=396050 $Y=64320
X9853 1 2 DECAP25JI3V $T=397040 24640 1 0 $X=396610 $Y=19520
X9854 1 2 DECAP25JI3V $T=397040 221760 1 0 $X=396610 $Y=216640
X9855 1 2 DECAP25JI3V $T=399280 194880 0 0 $X=398850 $Y=194240
X9856 1 2 DECAP25JI3V $T=400400 105280 0 0 $X=399970 $Y=104640
X9857 1 2 DECAP25JI3V $T=400400 123200 1 0 $X=399970 $Y=118080
X9858 1 2 DECAP25JI3V $T=400400 194880 1 0 $X=399970 $Y=189760
X9859 1 2 DECAP25JI3V $T=400400 212800 0 0 $X=399970 $Y=212160
X9860 1 2 DECAP25JI3V $T=401520 176960 1 0 $X=401090 $Y=171840
X9861 1 2 DECAP25JI3V $T=402640 185920 0 0 $X=402210 $Y=185280
X9862 1 2 DECAP25JI3V $T=403200 123200 0 0 $X=402770 $Y=122560
X9863 1 2 DECAP25JI3V $T=407120 42560 1 0 $X=406690 $Y=37440
X9864 1 2 DECAP25JI3V $T=407120 42560 0 0 $X=406690 $Y=41920
X9865 1 2 DECAP25JI3V $T=407120 51520 1 0 $X=406690 $Y=46400
X9866 1 2 DECAP25JI3V $T=407120 51520 0 0 $X=406690 $Y=50880
X9867 1 2 DECAP25JI3V $T=407120 60480 1 0 $X=406690 $Y=55360
X9868 1 2 DECAP25JI3V $T=407120 60480 0 0 $X=406690 $Y=59840
X9869 1 2 DECAP25JI3V $T=407120 69440 0 0 $X=406690 $Y=68800
X9870 1 2 DECAP25JI3V $T=407120 132160 1 0 $X=406690 $Y=127040
X9871 1 2 DECAP25JI3V $T=407120 159040 0 0 $X=406690 $Y=158400
X9872 1 2 DECAP25JI3V $T=407120 168000 1 0 $X=406690 $Y=162880
X9873 1 2 DECAP25JI3V $T=407120 168000 0 0 $X=406690 $Y=167360
X9874 1 2 DECAP25JI3V $T=408240 24640 0 0 $X=407810 $Y=24000
X9875 1 2 DECAP25JI3V $T=408240 159040 1 0 $X=407810 $Y=153920
X9876 1 2 DECAP25JI3V $T=411040 24640 1 0 $X=410610 $Y=19520
X9877 1 2 DECAP25JI3V $T=411040 221760 1 0 $X=410610 $Y=216640
X9878 1 2 DECAP10JI3V $T=20160 60480 0 0 $X=19730 $Y=59840
X9879 1 2 DECAP10JI3V $T=20160 69440 1 0 $X=19730 $Y=64320
X9880 1 2 DECAP10JI3V $T=20160 87360 1 0 $X=19730 $Y=82240
X9881 1 2 DECAP10JI3V $T=20160 96320 1 0 $X=19730 $Y=91200
X9882 1 2 DECAP10JI3V $T=20160 168000 0 0 $X=19730 $Y=167360
X9883 1 2 DECAP10JI3V $T=20160 212800 1 0 $X=19730 $Y=207680
X9884 1 2 DECAP10JI3V $T=24080 114240 0 0 $X=23650 $Y=113600
X9885 1 2 DECAP10JI3V $T=39200 141120 0 0 $X=38770 $Y=140480
X9886 1 2 DECAP10JI3V $T=48160 24640 1 0 $X=47730 $Y=19520
X9887 1 2 DECAP10JI3V $T=48160 87360 0 0 $X=47730 $Y=86720
X9888 1 2 DECAP10JI3V $T=48160 221760 1 0 $X=47730 $Y=216640
X9889 1 2 DECAP10JI3V $T=69440 78400 0 180 $X=63410 $Y=73280
X9890 1 2 DECAP10JI3V $T=68320 159040 0 0 $X=67890 $Y=158400
X9891 1 2 DECAP10JI3V $T=100800 176960 1 0 $X=100370 $Y=171840
X9892 1 2 DECAP10JI3V $T=104720 24640 0 0 $X=104290 $Y=24000
X9893 1 2 DECAP10JI3V $T=133280 176960 1 0 $X=132850 $Y=171840
X9894 1 2 DECAP10JI3V $T=148400 96320 1 0 $X=147970 $Y=91200
X9895 1 2 DECAP10JI3V $T=148400 141120 1 0 $X=147970 $Y=136000
X9896 1 2 DECAP10JI3V $T=197680 123200 0 0 $X=197250 $Y=122560
X9897 1 2 DECAP10JI3V $T=197680 132160 0 0 $X=197250 $Y=131520
X9898 1 2 DECAP10JI3V $T=205520 96320 0 0 $X=205090 $Y=95680
X9899 1 2 DECAP10JI3V $T=210000 123200 1 0 $X=209570 $Y=118080
X9900 1 2 DECAP10JI3V $T=210000 159040 1 0 $X=209570 $Y=153920
X9901 1 2 DECAP10JI3V $T=212800 24640 1 0 $X=212370 $Y=19520
X9902 1 2 DECAP10JI3V $T=213360 33600 1 0 $X=212930 $Y=28480
X9903 1 2 DECAP10JI3V $T=226240 105280 1 0 $X=225810 $Y=100160
X9904 1 2 DECAP10JI3V $T=239120 159040 0 0 $X=238690 $Y=158400
X9905 1 2 DECAP10JI3V $T=240240 96320 0 0 $X=239810 $Y=95680
X9906 1 2 DECAP10JI3V $T=246960 141120 1 0 $X=246530 $Y=136000
X9907 1 2 DECAP10JI3V $T=310240 141120 1 0 $X=309810 $Y=136000
X9908 1 2 DECAP10JI3V $T=315280 69440 0 0 $X=314850 $Y=68800
X9909 1 2 DECAP10JI3V $T=315280 87360 1 0 $X=314850 $Y=82240
X9910 1 2 DECAP10JI3V $T=316400 24640 1 0 $X=315970 $Y=19520
X9911 1 2 DECAP10JI3V $T=317520 159040 1 0 $X=317090 $Y=153920
X9912 1 2 DECAP10JI3V $T=317520 194880 0 0 $X=317090 $Y=194240
X9913 1 2 DECAP10JI3V $T=317520 203840 0 0 $X=317090 $Y=203200
X9914 1 2 DECAP10JI3V $T=318080 24640 0 0 $X=317650 $Y=24000
X9915 1 2 DECAP10JI3V $T=338800 159040 0 0 $X=338370 $Y=158400
X9916 1 2 DECAP10JI3V $T=351680 105280 1 0 $X=351250 $Y=100160
X9917 1 2 DECAP10JI3V $T=353360 96320 0 0 $X=352930 $Y=95680
X9918 1 2 DECAP10JI3V $T=403760 150080 1 0 $X=403330 $Y=144960
X9919 1 2 DECAP10JI3V $T=407680 33600 0 0 $X=407250 $Y=32960
X9920 1 2 DECAP10JI3V $T=415520 176960 1 0 $X=415090 $Y=171840
X9921 1 2 DECAP7JI3V $T=20160 33600 0 0 $X=19730 $Y=32960
X9922 1 2 DECAP7JI3V $T=20160 42560 1 0 $X=19730 $Y=37440
X9923 1 2 DECAP7JI3V $T=20160 51520 0 0 $X=19730 $Y=50880
X9924 1 2 DECAP7JI3V $T=20160 78400 1 0 $X=19730 $Y=73280
X9925 1 2 DECAP7JI3V $T=20160 78400 0 0 $X=19730 $Y=77760
X9926 1 2 DECAP7JI3V $T=20160 105280 1 0 $X=19730 $Y=100160
X9927 1 2 DECAP7JI3V $T=20160 105280 0 0 $X=19730 $Y=104640
X9928 1 2 DECAP7JI3V $T=20160 114240 1 0 $X=19730 $Y=109120
X9929 1 2 DECAP7JI3V $T=20160 114240 0 0 $X=19730 $Y=113600
X9930 1 2 DECAP7JI3V $T=20160 123200 0 0 $X=19730 $Y=122560
X9931 1 2 DECAP7JI3V $T=20160 141120 1 0 $X=19730 $Y=136000
X9932 1 2 DECAP7JI3V $T=20160 141120 0 0 $X=19730 $Y=140480
X9933 1 2 DECAP7JI3V $T=20160 159040 0 0 $X=19730 $Y=158400
X9934 1 2 DECAP7JI3V $T=20160 185920 1 0 $X=19730 $Y=180800
X9935 1 2 DECAP7JI3V $T=20160 185920 0 0 $X=19730 $Y=185280
X9936 1 2 DECAP7JI3V $T=20160 194880 0 0 $X=19730 $Y=194240
X9937 1 2 DECAP7JI3V $T=20160 203840 1 0 $X=19730 $Y=198720
X9938 1 2 DECAP7JI3V $T=24080 78400 0 0 $X=23650 $Y=77760
X9939 1 2 DECAP7JI3V $T=24080 159040 0 0 $X=23650 $Y=158400
X9940 1 2 DECAP7JI3V $T=24080 203840 1 0 $X=23650 $Y=198720
X9941 1 2 DECAP7JI3V $T=28000 203840 1 0 $X=27570 $Y=198720
X9942 1 2 DECAP7JI3V $T=31920 203840 1 0 $X=31490 $Y=198720
X9943 1 2 DECAP7JI3V $T=34160 24640 0 0 $X=33730 $Y=24000
X9944 1 2 DECAP7JI3V $T=34160 168000 1 0 $X=33730 $Y=162880
X9945 1 2 DECAP7JI3V $T=34720 114240 0 0 $X=34290 $Y=113600
X9946 1 2 DECAP7JI3V $T=34720 123200 1 0 $X=34290 $Y=118080
X9947 1 2 DECAP7JI3V $T=38080 24640 0 0 $X=37650 $Y=24000
X9948 1 2 DECAP7JI3V $T=38080 168000 1 0 $X=37650 $Y=162880
X9949 1 2 DECAP7JI3V $T=38640 123200 1 0 $X=38210 $Y=118080
X9950 1 2 DECAP7JI3V $T=42000 24640 0 0 $X=41570 $Y=24000
X9951 1 2 DECAP7JI3V $T=42000 168000 1 0 $X=41570 $Y=162880
X9952 1 2 DECAP7JI3V $T=43120 42560 0 0 $X=42690 $Y=41920
X9953 1 2 DECAP7JI3V $T=43120 78400 0 0 $X=42690 $Y=77760
X9954 1 2 DECAP7JI3V $T=43680 123200 1 0 $X=43250 $Y=118080
X9955 1 2 DECAP7JI3V $T=45920 24640 0 0 $X=45490 $Y=24000
X9956 1 2 DECAP7JI3V $T=49280 159040 0 0 $X=48850 $Y=158400
X9957 1 2 DECAP7JI3V $T=53760 24640 1 0 $X=53330 $Y=19520
X9958 1 2 DECAP7JI3V $T=53760 221760 1 0 $X=53330 $Y=216640
X9959 1 2 DECAP7JI3V $T=57680 24640 1 0 $X=57250 $Y=19520
X9960 1 2 DECAP7JI3V $T=57680 221760 1 0 $X=57250 $Y=216640
X9961 1 2 DECAP7JI3V $T=62720 150080 0 0 $X=62290 $Y=149440
X9962 1 2 DECAP7JI3V $T=64400 176960 1 0 $X=63970 $Y=171840
X9963 1 2 DECAP7JI3V $T=69440 78400 1 0 $X=69010 $Y=73280
X9964 1 2 DECAP7JI3V $T=77280 60480 0 0 $X=76850 $Y=59840
X9965 1 2 DECAP7JI3V $T=92960 33600 0 180 $X=88610 $Y=28480
X9966 1 2 DECAP7JI3V $T=94640 87360 1 0 $X=94210 $Y=82240
X9967 1 2 DECAP7JI3V $T=101360 60480 1 0 $X=100930 $Y=55360
X9968 1 2 DECAP7JI3V $T=101360 60480 0 0 $X=100930 $Y=59840
X9969 1 2 DECAP7JI3V $T=101360 69440 1 0 $X=100930 $Y=64320
X9970 1 2 DECAP7JI3V $T=101360 69440 0 0 $X=100930 $Y=68800
X9971 1 2 DECAP7JI3V $T=101360 78400 1 0 $X=100930 $Y=73280
X9972 1 2 DECAP7JI3V $T=101360 168000 0 0 $X=100930 $Y=167360
X9973 1 2 DECAP7JI3V $T=103040 105280 0 0 $X=102610 $Y=104640
X9974 1 2 DECAP7JI3V $T=105280 24640 1 0 $X=104850 $Y=19520
X9975 1 2 DECAP7JI3V $T=105280 42560 0 0 $X=104850 $Y=41920
X9976 1 2 DECAP7JI3V $T=105280 51520 0 0 $X=104850 $Y=50880
X9977 1 2 DECAP7JI3V $T=105280 60480 1 0 $X=104850 $Y=55360
X9978 1 2 DECAP7JI3V $T=105280 60480 0 0 $X=104850 $Y=59840
X9979 1 2 DECAP7JI3V $T=105280 69440 1 0 $X=104850 $Y=64320
X9980 1 2 DECAP7JI3V $T=105280 69440 0 0 $X=104850 $Y=68800
X9981 1 2 DECAP7JI3V $T=105280 78400 1 0 $X=104850 $Y=73280
X9982 1 2 DECAP7JI3V $T=105280 87360 1 0 $X=104850 $Y=82240
X9983 1 2 DECAP7JI3V $T=105280 132160 1 0 $X=104850 $Y=127040
X9984 1 2 DECAP7JI3V $T=105280 132160 0 0 $X=104850 $Y=131520
X9985 1 2 DECAP7JI3V $T=105280 141120 1 0 $X=104850 $Y=136000
X9986 1 2 DECAP7JI3V $T=105280 141120 0 0 $X=104850 $Y=140480
X9987 1 2 DECAP7JI3V $T=105280 150080 1 0 $X=104850 $Y=144960
X9988 1 2 DECAP7JI3V $T=105280 194880 0 0 $X=104850 $Y=194240
X9989 1 2 DECAP7JI3V $T=106400 176960 1 0 $X=105970 $Y=171840
X9990 1 2 DECAP7JI3V $T=106960 105280 0 0 $X=106530 $Y=104640
X9991 1 2 DECAP7JI3V $T=109200 24640 1 0 $X=108770 $Y=19520
X9992 1 2 DECAP7JI3V $T=109200 60480 1 0 $X=108770 $Y=55360
X9993 1 2 DECAP7JI3V $T=109200 60480 0 0 $X=108770 $Y=59840
X9994 1 2 DECAP7JI3V $T=109200 69440 1 0 $X=108770 $Y=64320
X9995 1 2 DECAP7JI3V $T=109200 69440 0 0 $X=108770 $Y=68800
X9996 1 2 DECAP7JI3V $T=109200 78400 1 0 $X=108770 $Y=73280
X9997 1 2 DECAP7JI3V $T=109200 87360 1 0 $X=108770 $Y=82240
X9998 1 2 DECAP7JI3V $T=109200 132160 1 0 $X=108770 $Y=127040
X9999 1 2 DECAP7JI3V $T=109200 132160 0 0 $X=108770 $Y=131520
X10000 1 2 DECAP7JI3V $T=109200 141120 1 0 $X=108770 $Y=136000
X10001 1 2 DECAP7JI3V $T=109200 141120 0 0 $X=108770 $Y=140480
X10002 1 2 DECAP7JI3V $T=109200 150080 1 0 $X=108770 $Y=144960
X10003 1 2 DECAP7JI3V $T=109200 159040 0 0 $X=108770 $Y=158400
X10004 1 2 DECAP7JI3V $T=109200 194880 0 0 $X=108770 $Y=194240
X10005 1 2 DECAP7JI3V $T=110320 176960 1 0 $X=109890 $Y=171840
X10006 1 2 DECAP7JI3V $T=114240 176960 1 0 $X=113810 $Y=171840
X10007 1 2 DECAP7JI3V $T=118720 78400 1 0 $X=118290 $Y=73280
X10008 1 2 DECAP7JI3V $T=118720 150080 0 0 $X=118290 $Y=149440
X10009 1 2 DECAP7JI3V $T=118720 212800 1 0 $X=118290 $Y=207680
X10010 1 2 DECAP7JI3V $T=118720 221760 1 0 $X=118290 $Y=216640
X10011 1 2 DECAP7JI3V $T=123200 168000 1 0 $X=122770 $Y=162880
X10012 1 2 DECAP7JI3V $T=123200 168000 0 0 $X=122770 $Y=167360
X10013 1 2 DECAP7JI3V $T=127120 212800 1 180 $X=122770 $Y=212160
X10014 1 2 DECAP7JI3V $T=127120 212800 0 0 $X=126690 $Y=212160
X10015 1 2 DECAP7JI3V $T=132720 33600 1 180 $X=128370 $Y=32960
X10016 1 2 DECAP7JI3V $T=131040 212800 0 0 $X=130610 $Y=212160
X10017 1 2 DECAP7JI3V $T=132720 185920 1 0 $X=132290 $Y=180800
X10018 1 2 DECAP7JI3V $T=133280 132160 0 0 $X=132850 $Y=131520
X10019 1 2 DECAP7JI3V $T=134960 212800 0 0 $X=134530 $Y=212160
X10020 1 2 DECAP7JI3V $T=149520 78400 0 0 $X=149090 $Y=77760
X10021 1 2 DECAP7JI3V $T=153440 78400 0 0 $X=153010 $Y=77760
X10022 1 2 DECAP7JI3V $T=154000 96320 1 0 $X=153570 $Y=91200
X10023 1 2 DECAP7JI3V $T=157360 78400 0 0 $X=156930 $Y=77760
X10024 1 2 DECAP7JI3V $T=157920 96320 1 0 $X=157490 $Y=91200
X10025 1 2 DECAP7JI3V $T=159040 123200 1 0 $X=158610 $Y=118080
X10026 1 2 DECAP7JI3V $T=161280 78400 0 0 $X=160850 $Y=77760
X10027 1 2 DECAP7JI3V $T=161840 96320 1 0 $X=161410 $Y=91200
X10028 1 2 DECAP7JI3V $T=162960 123200 1 0 $X=162530 $Y=118080
X10029 1 2 DECAP7JI3V $T=167440 105280 1 0 $X=167010 $Y=100160
X10030 1 2 DECAP7JI3V $T=174160 33600 0 0 $X=173730 $Y=32960
X10031 1 2 DECAP7JI3V $T=175840 141120 0 0 $X=175410 $Y=140480
X10032 1 2 DECAP7JI3V $T=179200 132160 1 0 $X=178770 $Y=127040
X10033 1 2 DECAP7JI3V $T=180320 105280 0 0 $X=179890 $Y=104640
X10034 1 2 DECAP7JI3V $T=182560 78400 1 0 $X=182130 $Y=73280
X10035 1 2 DECAP7JI3V $T=184240 33600 1 0 $X=183810 $Y=28480
X10036 1 2 DECAP7JI3V $T=184240 60480 1 0 $X=183810 $Y=55360
X10037 1 2 DECAP7JI3V $T=184240 105280 0 0 $X=183810 $Y=104640
X10038 1 2 DECAP7JI3V $T=185920 87360 1 0 $X=185490 $Y=82240
X10039 1 2 DECAP7JI3V $T=185920 132160 1 0 $X=185490 $Y=127040
X10040 1 2 DECAP7JI3V $T=190400 78400 0 180 $X=186050 $Y=73280
X10041 1 2 DECAP7JI3V $T=189840 87360 1 0 $X=189410 $Y=82240
X10042 1 2 DECAP7JI3V $T=194880 60480 0 0 $X=194450 $Y=59840
X10043 1 2 DECAP7JI3V $T=203280 123200 0 0 $X=202850 $Y=122560
X10044 1 2 DECAP7JI3V $T=203280 132160 0 0 $X=202850 $Y=131520
X10045 1 2 DECAP7JI3V $T=206080 168000 1 0 $X=205650 $Y=162880
X10046 1 2 DECAP7JI3V $T=206080 168000 0 0 $X=205650 $Y=167360
X10047 1 2 DECAP7JI3V $T=206080 176960 1 0 $X=205650 $Y=171840
X10048 1 2 DECAP7JI3V $T=207200 123200 0 0 $X=206770 $Y=122560
X10049 1 2 DECAP7JI3V $T=207200 132160 0 0 $X=206770 $Y=131520
X10050 1 2 DECAP7JI3V $T=207200 150080 0 0 $X=206770 $Y=149440
X10051 1 2 DECAP7JI3V $T=208320 105280 0 0 $X=207890 $Y=104640
X10052 1 2 DECAP7JI3V $T=210000 168000 1 0 $X=209570 $Y=162880
X10053 1 2 DECAP7JI3V $T=210000 168000 0 0 $X=209570 $Y=167360
X10054 1 2 DECAP7JI3V $T=210000 176960 1 0 $X=209570 $Y=171840
X10055 1 2 DECAP7JI3V $T=211120 96320 0 0 $X=210690 $Y=95680
X10056 1 2 DECAP7JI3V $T=211120 123200 0 0 $X=210690 $Y=122560
X10057 1 2 DECAP7JI3V $T=211120 132160 1 0 $X=210690 $Y=127040
X10058 1 2 DECAP7JI3V $T=211120 132160 0 0 $X=210690 $Y=131520
X10059 1 2 DECAP7JI3V $T=211120 150080 0 0 $X=210690 $Y=149440
X10060 1 2 DECAP7JI3V $T=212240 105280 0 0 $X=211810 $Y=104640
X10061 1 2 DECAP7JI3V $T=213920 114240 0 0 $X=213490 $Y=113600
X10062 1 2 DECAP7JI3V $T=215040 96320 0 0 $X=214610 $Y=95680
X10063 1 2 DECAP7JI3V $T=215040 123200 0 0 $X=214610 $Y=122560
X10064 1 2 DECAP7JI3V $T=215040 132160 1 0 $X=214610 $Y=127040
X10065 1 2 DECAP7JI3V $T=215040 132160 0 0 $X=214610 $Y=131520
X10066 1 2 DECAP7JI3V $T=215040 141120 1 0 $X=214610 $Y=136000
X10067 1 2 DECAP7JI3V $T=215040 150080 0 0 $X=214610 $Y=149440
X10068 1 2 DECAP7JI3V $T=215040 159040 0 0 $X=214610 $Y=158400
X10069 1 2 DECAP7JI3V $T=215040 176960 0 0 $X=214610 $Y=176320
X10070 1 2 DECAP7JI3V $T=218960 141120 1 0 $X=218530 $Y=136000
X10071 1 2 DECAP7JI3V $T=236320 42560 1 0 $X=235890 $Y=37440
X10072 1 2 DECAP7JI3V $T=243600 87360 1 0 $X=243170 $Y=82240
X10073 1 2 DECAP7JI3V $T=254800 168000 1 180 $X=250450 $Y=167360
X10074 1 2 DECAP7JI3V $T=253680 141120 1 0 $X=253250 $Y=136000
X10075 1 2 DECAP7JI3V $T=261520 141120 0 180 $X=257170 $Y=136000
X10076 1 2 DECAP7JI3V $T=260400 87360 0 0 $X=259970 $Y=86720
X10077 1 2 DECAP7JI3V $T=260400 123200 1 0 $X=259970 $Y=118080
X10078 1 2 DECAP7JI3V $T=260400 123200 0 0 $X=259970 $Y=122560
X10079 1 2 DECAP7JI3V $T=260960 132160 1 0 $X=260530 $Y=127040
X10080 1 2 DECAP7JI3V $T=264320 87360 0 0 $X=263890 $Y=86720
X10081 1 2 DECAP7JI3V $T=268240 87360 0 0 $X=267810 $Y=86720
X10082 1 2 DECAP7JI3V $T=277200 176960 0 0 $X=276770 $Y=176320
X10083 1 2 DECAP7JI3V $T=278880 78400 0 0 $X=278450 $Y=77760
X10084 1 2 DECAP7JI3V $T=282240 105280 1 0 $X=281810 $Y=100160
X10085 1 2 DECAP7JI3V $T=282240 114240 1 0 $X=281810 $Y=109120
X10086 1 2 DECAP7JI3V $T=282800 78400 0 0 $X=282370 $Y=77760
X10087 1 2 DECAP7JI3V $T=284480 123200 0 0 $X=284050 $Y=122560
X10088 1 2 DECAP7JI3V $T=285040 132160 0 0 $X=284610 $Y=131520
X10089 1 2 DECAP7JI3V $T=286160 105280 1 0 $X=285730 $Y=100160
X10090 1 2 DECAP7JI3V $T=290080 105280 1 0 $X=289650 $Y=100160
X10091 1 2 DECAP7JI3V $T=290640 96320 1 0 $X=290210 $Y=91200
X10092 1 2 DECAP7JI3V $T=293440 87360 0 0 $X=293010 $Y=86720
X10093 1 2 DECAP7JI3V $T=297360 87360 0 0 $X=296930 $Y=86720
X10094 1 2 DECAP7JI3V $T=305760 42560 0 0 $X=305330 $Y=41920
X10095 1 2 DECAP7JI3V $T=306880 42560 1 0 $X=306450 $Y=37440
X10096 1 2 DECAP7JI3V $T=307440 150080 1 0 $X=307010 $Y=144960
X10097 1 2 DECAP7JI3V $T=309120 78400 1 0 $X=308690 $Y=73280
X10098 1 2 DECAP7JI3V $T=309120 96320 0 0 $X=308690 $Y=95680
X10099 1 2 DECAP7JI3V $T=309120 105280 1 0 $X=308690 $Y=100160
X10100 1 2 DECAP7JI3V $T=309120 114240 1 0 $X=308690 $Y=109120
X10101 1 2 DECAP7JI3V $T=309120 141120 0 0 $X=308690 $Y=140480
X10102 1 2 DECAP7JI3V $T=313040 78400 1 0 $X=312610 $Y=73280
X10103 1 2 DECAP7JI3V $T=313040 96320 0 0 $X=312610 $Y=95680
X10104 1 2 DECAP7JI3V $T=313040 105280 1 0 $X=312610 $Y=100160
X10105 1 2 DECAP7JI3V $T=313040 114240 1 0 $X=312610 $Y=109120
X10106 1 2 DECAP7JI3V $T=313040 141120 0 0 $X=312610 $Y=140480
X10107 1 2 DECAP7JI3V $T=315840 141120 1 0 $X=315410 $Y=136000
X10108 1 2 DECAP7JI3V $T=315840 159040 0 0 $X=315410 $Y=158400
X10109 1 2 DECAP7JI3V $T=315840 168000 1 0 $X=315410 $Y=162880
X10110 1 2 DECAP7JI3V $T=316960 78400 1 0 $X=316530 $Y=73280
X10111 1 2 DECAP7JI3V $T=316960 123200 1 0 $X=316530 $Y=118080
X10112 1 2 DECAP7JI3V $T=316960 132160 1 0 $X=316530 $Y=127040
X10113 1 2 DECAP7JI3V $T=316960 150080 1 0 $X=316530 $Y=144960
X10114 1 2 DECAP7JI3V $T=318080 87360 0 0 $X=317650 $Y=86720
X10115 1 2 DECAP7JI3V $T=318080 123200 0 0 $X=317650 $Y=122560
X10116 1 2 DECAP7JI3V $T=319200 42560 0 0 $X=318770 $Y=41920
X10117 1 2 DECAP7JI3V $T=320880 69440 0 0 $X=320450 $Y=68800
X10118 1 2 DECAP7JI3V $T=320880 78400 1 0 $X=320450 $Y=73280
X10119 1 2 DECAP7JI3V $T=320880 87360 1 0 $X=320450 $Y=82240
X10120 1 2 DECAP7JI3V $T=320880 123200 1 0 $X=320450 $Y=118080
X10121 1 2 DECAP7JI3V $T=320880 132160 1 0 $X=320450 $Y=127040
X10122 1 2 DECAP7JI3V $T=320880 150080 1 0 $X=320450 $Y=144960
X10123 1 2 DECAP7JI3V $T=322000 212800 1 0 $X=321570 $Y=207680
X10124 1 2 DECAP7JI3V $T=329840 132160 0 0 $X=329410 $Y=131520
X10125 1 2 DECAP7JI3V $T=330400 78400 0 0 $X=329970 $Y=77760
X10126 1 2 DECAP7JI3V $T=330400 105280 0 0 $X=329970 $Y=104640
X10127 1 2 DECAP7JI3V $T=334320 78400 0 0 $X=333890 $Y=77760
X10128 1 2 DECAP7JI3V $T=344960 114240 0 0 $X=344530 $Y=113600
X10129 1 2 DECAP7JI3V $T=348880 114240 0 0 $X=348450 $Y=113600
X10130 1 2 DECAP7JI3V $T=352800 114240 0 0 $X=352370 $Y=113600
X10131 1 2 DECAP7JI3V $T=352800 141120 0 0 $X=352370 $Y=140480
X10132 1 2 DECAP7JI3V $T=356720 114240 1 0 $X=356290 $Y=109120
X10133 1 2 DECAP7JI3V $T=356720 114240 0 0 $X=356290 $Y=113600
X10134 1 2 DECAP7JI3V $T=356720 141120 0 0 $X=356290 $Y=140480
X10135 1 2 DECAP7JI3V $T=357280 42560 0 0 $X=356850 $Y=41920
X10136 1 2 DECAP7JI3V $T=357280 51520 1 0 $X=356850 $Y=46400
X10137 1 2 DECAP7JI3V $T=358400 96320 1 0 $X=357970 $Y=91200
X10138 1 2 DECAP7JI3V $T=358960 60480 1 0 $X=358530 $Y=55360
X10139 1 2 DECAP7JI3V $T=359520 78400 0 0 $X=359090 $Y=77760
X10140 1 2 DECAP7JI3V $T=360080 69440 0 0 $X=359650 $Y=68800
X10141 1 2 DECAP7JI3V $T=406560 78400 0 0 $X=406130 $Y=77760
X10142 1 2 DECAP7JI3V $T=406560 87360 0 0 $X=406130 $Y=86720
X10143 1 2 DECAP7JI3V $T=406560 96320 1 0 $X=406130 $Y=91200
X10144 1 2 DECAP7JI3V $T=406560 150080 0 0 $X=406130 $Y=149440
X10145 1 2 DECAP7JI3V $T=409360 78400 1 0 $X=408930 $Y=73280
X10146 1 2 DECAP7JI3V $T=409360 87360 1 0 $X=408930 $Y=82240
X10147 1 2 DECAP7JI3V $T=409360 150080 1 0 $X=408930 $Y=144960
X10148 1 2 DECAP7JI3V $T=409360 203840 1 0 $X=408930 $Y=198720
X10149 1 2 DECAP7JI3V $T=409360 212800 1 0 $X=408930 $Y=207680
X10150 1 2 DECAP7JI3V $T=410480 69440 1 0 $X=410050 $Y=64320
X10151 1 2 DECAP7JI3V $T=410480 78400 0 0 $X=410050 $Y=77760
X10152 1 2 DECAP7JI3V $T=410480 87360 0 0 $X=410050 $Y=86720
X10153 1 2 DECAP7JI3V $T=410480 96320 1 0 $X=410050 $Y=91200
X10154 1 2 DECAP7JI3V $T=410480 150080 0 0 $X=410050 $Y=149440
X10155 1 2 DECAP7JI3V $T=410480 185920 1 0 $X=410050 $Y=180800
X10156 1 2 DECAP7JI3V $T=413280 33600 0 0 $X=412850 $Y=32960
X10157 1 2 DECAP7JI3V $T=413280 78400 1 0 $X=412850 $Y=73280
X10158 1 2 DECAP7JI3V $T=413280 87360 1 0 $X=412850 $Y=82240
X10159 1 2 DECAP7JI3V $T=413280 150080 1 0 $X=412850 $Y=144960
X10160 1 2 DECAP7JI3V $T=413280 194880 0 0 $X=412850 $Y=194240
X10161 1 2 DECAP7JI3V $T=413280 203840 1 0 $X=412850 $Y=198720
X10162 1 2 DECAP7JI3V $T=413280 203840 0 0 $X=412850 $Y=203200
X10163 1 2 DECAP7JI3V $T=413280 212800 1 0 $X=412850 $Y=207680
X10164 1 2 DECAP7JI3V $T=414400 69440 1 0 $X=413970 $Y=64320
X10165 1 2 DECAP7JI3V $T=414400 78400 0 0 $X=413970 $Y=77760
X10166 1 2 DECAP7JI3V $T=414400 87360 0 0 $X=413970 $Y=86720
X10167 1 2 DECAP7JI3V $T=414400 96320 1 0 $X=413970 $Y=91200
X10168 1 2 DECAP7JI3V $T=414400 105280 0 0 $X=413970 $Y=104640
X10169 1 2 DECAP7JI3V $T=414400 123200 1 0 $X=413970 $Y=118080
X10170 1 2 DECAP7JI3V $T=414400 150080 0 0 $X=413970 $Y=149440
X10171 1 2 DECAP7JI3V $T=414400 176960 0 0 $X=413970 $Y=176320
X10172 1 2 DECAP7JI3V $T=414400 185920 1 0 $X=413970 $Y=180800
X10173 1 2 DECAP7JI3V $T=414400 194880 1 0 $X=413970 $Y=189760
X10174 1 2 DECAP7JI3V $T=414400 212800 0 0 $X=413970 $Y=212160
X10175 1 2 DECAP7JI3V $T=417200 33600 1 0 $X=416770 $Y=28480
X10176 1 2 DECAP7JI3V $T=417200 33600 0 0 $X=416770 $Y=32960
X10177 1 2 DECAP7JI3V $T=417200 78400 1 0 $X=416770 $Y=73280
X10178 1 2 DECAP7JI3V $T=417200 87360 1 0 $X=416770 $Y=82240
X10179 1 2 DECAP7JI3V $T=417200 114240 1 0 $X=416770 $Y=109120
X10180 1 2 DECAP7JI3V $T=417200 123200 0 0 $X=416770 $Y=122560
X10181 1 2 DECAP7JI3V $T=417200 141120 0 0 $X=416770 $Y=140480
X10182 1 2 DECAP7JI3V $T=417200 150080 1 0 $X=416770 $Y=144960
X10183 1 2 DECAP7JI3V $T=417200 194880 0 0 $X=416770 $Y=194240
X10184 1 2 DECAP7JI3V $T=417200 203840 1 0 $X=416770 $Y=198720
X10185 1 2 DECAP7JI3V $T=417200 203840 0 0 $X=416770 $Y=203200
X10186 1 2 DECAP7JI3V $T=417200 212800 1 0 $X=416770 $Y=207680
X10187 1 2 DECAP7JI3V $T=418320 69440 1 0 $X=417890 $Y=64320
X10188 1 2 DECAP7JI3V $T=418320 78400 0 0 $X=417890 $Y=77760
X10189 1 2 DECAP7JI3V $T=418320 87360 0 0 $X=417890 $Y=86720
X10190 1 2 DECAP7JI3V $T=418320 96320 1 0 $X=417890 $Y=91200
X10191 1 2 DECAP7JI3V $T=418320 96320 0 0 $X=417890 $Y=95680
X10192 1 2 DECAP7JI3V $T=418320 105280 1 0 $X=417890 $Y=100160
X10193 1 2 DECAP7JI3V $T=418320 105280 0 0 $X=417890 $Y=104640
X10194 1 2 DECAP7JI3V $T=418320 114240 0 0 $X=417890 $Y=113600
X10195 1 2 DECAP7JI3V $T=418320 123200 1 0 $X=417890 $Y=118080
X10196 1 2 DECAP7JI3V $T=418320 132160 0 0 $X=417890 $Y=131520
X10197 1 2 DECAP7JI3V $T=418320 141120 1 0 $X=417890 $Y=136000
X10198 1 2 DECAP7JI3V $T=418320 150080 0 0 $X=417890 $Y=149440
X10199 1 2 DECAP7JI3V $T=418320 176960 0 0 $X=417890 $Y=176320
X10200 1 2 DECAP7JI3V $T=418320 185920 1 0 $X=417890 $Y=180800
X10201 1 2 DECAP7JI3V $T=418320 194880 1 0 $X=417890 $Y=189760
X10202 1 2 DECAP7JI3V $T=418320 212800 0 0 $X=417890 $Y=212160
X10203 1 2 DECAP7JI3V $T=421120 33600 1 0 $X=420690 $Y=28480
X10204 1 2 DECAP7JI3V $T=421120 33600 0 0 $X=420690 $Y=32960
X10205 1 2 DECAP7JI3V $T=421120 42560 1 0 $X=420690 $Y=37440
X10206 1 2 DECAP7JI3V $T=421120 42560 0 0 $X=420690 $Y=41920
X10207 1 2 DECAP7JI3V $T=421120 51520 1 0 $X=420690 $Y=46400
X10208 1 2 DECAP7JI3V $T=421120 51520 0 0 $X=420690 $Y=50880
X10209 1 2 DECAP7JI3V $T=421120 60480 1 0 $X=420690 $Y=55360
X10210 1 2 DECAP7JI3V $T=421120 60480 0 0 $X=420690 $Y=59840
X10211 1 2 DECAP7JI3V $T=421120 69440 0 0 $X=420690 $Y=68800
X10212 1 2 DECAP7JI3V $T=421120 78400 1 0 $X=420690 $Y=73280
X10213 1 2 DECAP7JI3V $T=421120 87360 1 0 $X=420690 $Y=82240
X10214 1 2 DECAP7JI3V $T=421120 114240 1 0 $X=420690 $Y=109120
X10215 1 2 DECAP7JI3V $T=421120 123200 0 0 $X=420690 $Y=122560
X10216 1 2 DECAP7JI3V $T=421120 132160 1 0 $X=420690 $Y=127040
X10217 1 2 DECAP7JI3V $T=421120 141120 0 0 $X=420690 $Y=140480
X10218 1 2 DECAP7JI3V $T=421120 150080 1 0 $X=420690 $Y=144960
X10219 1 2 DECAP7JI3V $T=421120 159040 0 0 $X=420690 $Y=158400
X10220 1 2 DECAP7JI3V $T=421120 168000 1 0 $X=420690 $Y=162880
X10221 1 2 DECAP7JI3V $T=421120 168000 0 0 $X=420690 $Y=167360
X10222 1 2 DECAP7JI3V $T=421120 176960 1 0 $X=420690 $Y=171840
X10223 1 2 DECAP7JI3V $T=421120 194880 0 0 $X=420690 $Y=194240
X10224 1 2 DECAP7JI3V $T=421120 203840 1 0 $X=420690 $Y=198720
X10225 1 2 DECAP7JI3V $T=421120 203840 0 0 $X=420690 $Y=203200
X10226 1 2 DECAP7JI3V $T=421120 212800 1 0 $X=420690 $Y=207680
X10227 1 2 DECAP5JI3V $T=20160 42560 0 0 $X=19730 $Y=41920
X10228 1 2 DECAP5JI3V $T=20160 51520 1 0 $X=19730 $Y=46400
X10229 1 2 DECAP5JI3V $T=20160 96320 0 0 $X=19730 $Y=95680
X10230 1 2 DECAP5JI3V $T=20160 132160 1 0 $X=19730 $Y=127040
X10231 1 2 DECAP5JI3V $T=20160 159040 1 0 $X=19730 $Y=153920
X10232 1 2 DECAP5JI3V $T=20160 176960 1 0 $X=19730 $Y=171840
X10233 1 2 DECAP5JI3V $T=30800 78400 1 180 $X=27570 $Y=77760
X10234 1 2 DECAP5JI3V $T=28560 203840 0 0 $X=28130 $Y=203200
X10235 1 2 DECAP5JI3V $T=34720 132160 1 0 $X=34290 $Y=127040
X10236 1 2 DECAP5JI3V $T=38640 203840 0 180 $X=35410 $Y=198720
X10237 1 2 DECAP5JI3V $T=39200 123200 0 0 $X=38770 $Y=122560
X10238 1 2 DECAP5JI3V $T=40880 96320 1 0 $X=40450 $Y=91200
X10239 1 2 DECAP5JI3V $T=42560 212800 0 0 $X=42130 $Y=212160
X10240 1 2 DECAP5JI3V $T=49840 24640 0 0 $X=49410 $Y=24000
X10241 1 2 DECAP5JI3V $T=57120 51520 0 0 $X=56690 $Y=50880
X10242 1 2 DECAP5JI3V $T=59360 60480 0 0 $X=58930 $Y=59840
X10243 1 2 DECAP5JI3V $T=59360 87360 1 0 $X=58930 $Y=82240
X10244 1 2 DECAP5JI3V $T=61040 33600 1 0 $X=60610 $Y=28480
X10245 1 2 DECAP5JI3V $T=66640 150080 0 0 $X=66210 $Y=149440
X10246 1 2 DECAP5JI3V $T=76720 60480 1 0 $X=76290 $Y=55360
X10247 1 2 DECAP5JI3V $T=78400 33600 0 0 $X=77970 $Y=32960
X10248 1 2 DECAP5JI3V $T=84000 105280 0 0 $X=83570 $Y=104640
X10249 1 2 DECAP5JI3V $T=105280 105280 1 0 $X=104850 $Y=100160
X10250 1 2 DECAP5JI3V $T=105280 168000 0 0 $X=104850 $Y=167360
X10251 1 2 DECAP5JI3V $T=105280 176960 0 0 $X=104850 $Y=176320
X10252 1 2 DECAP5JI3V $T=105280 212800 0 0 $X=104850 $Y=212160
X10253 1 2 DECAP5JI3V $T=108640 150080 0 0 $X=108210 $Y=149440
X10254 1 2 DECAP5JI3V $T=108640 159040 1 0 $X=108210 $Y=153920
X10255 1 2 DECAP5JI3V $T=110320 96320 0 0 $X=109890 $Y=95680
X10256 1 2 DECAP5JI3V $T=110320 203840 1 0 $X=109890 $Y=198720
X10257 1 2 DECAP5JI3V $T=113120 123200 1 0 $X=112690 $Y=118080
X10258 1 2 DECAP5JI3V $T=113120 159040 0 0 $X=112690 $Y=158400
X10259 1 2 DECAP5JI3V $T=122640 78400 1 0 $X=122210 $Y=73280
X10260 1 2 DECAP5JI3V $T=122640 150080 0 0 $X=122210 $Y=149440
X10261 1 2 DECAP5JI3V $T=133280 114240 0 0 $X=132850 $Y=113600
X10262 1 2 DECAP5JI3V $T=143360 212800 1 0 $X=142930 $Y=207680
X10263 1 2 DECAP5JI3V $T=156240 132160 1 0 $X=155810 $Y=127040
X10264 1 2 DECAP5JI3V $T=164080 87360 1 0 $X=163650 $Y=82240
X10265 1 2 DECAP5JI3V $T=166880 123200 1 0 $X=166450 $Y=118080
X10266 1 2 DECAP5JI3V $T=168560 96320 0 0 $X=168130 $Y=95680
X10267 1 2 DECAP5JI3V $T=179760 141120 0 0 $X=179330 $Y=140480
X10268 1 2 DECAP5JI3V $T=188160 150080 1 0 $X=187730 $Y=144960
X10269 1 2 DECAP5JI3V $T=190960 168000 1 180 $X=187730 $Y=167360
X10270 1 2 DECAP5JI3V $T=188160 176960 1 0 $X=187730 $Y=171840
X10271 1 2 DECAP5JI3V $T=211120 185920 1 0 $X=210690 $Y=180800
X10272 1 2 DECAP5JI3V $T=211120 212800 1 0 $X=210690 $Y=207680
X10273 1 2 DECAP5JI3V $T=211680 42560 0 0 $X=211250 $Y=41920
X10274 1 2 DECAP5JI3V $T=211680 51520 1 0 $X=211250 $Y=46400
X10275 1 2 DECAP5JI3V $T=211680 60480 1 0 $X=211250 $Y=55360
X10276 1 2 DECAP5JI3V $T=211680 69440 0 0 $X=211250 $Y=68800
X10277 1 2 DECAP5JI3V $T=211680 78400 0 0 $X=211250 $Y=77760
X10278 1 2 DECAP5JI3V $T=214480 87360 0 0 $X=214050 $Y=86720
X10279 1 2 DECAP5JI3V $T=214480 150080 1 0 $X=214050 $Y=144960
X10280 1 2 DECAP5JI3V $T=215040 212800 0 0 $X=214610 $Y=212160
X10281 1 2 DECAP5JI3V $T=216160 96320 1 0 $X=215730 $Y=91200
X10282 1 2 DECAP5JI3V $T=216160 105280 0 0 $X=215730 $Y=104640
X10283 1 2 DECAP5JI3V $T=229600 42560 0 0 $X=229170 $Y=41920
X10284 1 2 DECAP5JI3V $T=232400 51520 0 180 $X=229170 $Y=46400
X10285 1 2 DECAP5JI3V $T=229600 60480 1 0 $X=229170 $Y=55360
X10286 1 2 DECAP5JI3V $T=230720 168000 1 0 $X=230290 $Y=162880
X10287 1 2 DECAP5JI3V $T=239120 141120 0 0 $X=238690 $Y=140480
X10288 1 2 DECAP5JI3V $T=247520 51520 0 0 $X=247090 $Y=50880
X10289 1 2 DECAP5JI3V $T=250320 60480 0 180 $X=247090 $Y=55360
X10290 1 2 DECAP5JI3V $T=261520 141120 1 0 $X=261090 $Y=136000
X10291 1 2 DECAP5JI3V $T=267680 96320 1 0 $X=267250 $Y=91200
X10292 1 2 DECAP5JI3V $T=269360 78400 1 0 $X=268930 $Y=73280
X10293 1 2 DECAP5JI3V $T=274400 114240 0 0 $X=273970 $Y=113600
X10294 1 2 DECAP5JI3V $T=284480 105280 0 0 $X=284050 $Y=104640
X10295 1 2 DECAP5JI3V $T=285600 123200 1 0 $X=285170 $Y=118080
X10296 1 2 DECAP5JI3V $T=286160 114240 1 0 $X=285730 $Y=109120
X10297 1 2 DECAP5JI3V $T=286160 141120 1 0 $X=285730 $Y=136000
X10298 1 2 DECAP5JI3V $T=289520 78400 1 180 $X=286290 $Y=77760
X10299 1 2 DECAP5JI3V $T=291200 96320 0 0 $X=290770 $Y=95680
X10300 1 2 DECAP5JI3V $T=301280 87360 0 0 $X=300850 $Y=86720
X10301 1 2 DECAP5JI3V $T=309120 194880 1 0 $X=308690 $Y=189760
X10302 1 2 DECAP5JI3V $T=316960 51520 0 0 $X=316530 $Y=50880
X10303 1 2 DECAP5JI3V $T=316960 60480 1 0 $X=316530 $Y=55360
X10304 1 2 DECAP5JI3V $T=316960 60480 0 0 $X=316530 $Y=59840
X10305 1 2 DECAP5JI3V $T=316960 69440 1 0 $X=316530 $Y=64320
X10306 1 2 DECAP5JI3V $T=316960 96320 0 0 $X=316530 $Y=95680
X10307 1 2 DECAP5JI3V $T=316960 105280 1 0 $X=316530 $Y=100160
X10308 1 2 DECAP5JI3V $T=316960 114240 1 0 $X=316530 $Y=109120
X10309 1 2 DECAP5JI3V $T=316960 141120 0 0 $X=316530 $Y=140480
X10310 1 2 DECAP5JI3V $T=316960 150080 0 0 $X=316530 $Y=149440
X10311 1 2 DECAP5JI3V $T=320320 105280 0 0 $X=319890 $Y=104640
X10312 1 2 DECAP5JI3V $T=322000 87360 0 0 $X=321570 $Y=86720
X10313 1 2 DECAP5JI3V $T=322000 114240 0 0 $X=321570 $Y=113600
X10314 1 2 DECAP5JI3V $T=322000 123200 0 0 $X=321570 $Y=122560
X10315 1 2 DECAP5JI3V $T=322000 212800 0 0 $X=321570 $Y=212160
X10316 1 2 DECAP5JI3V $T=323120 132160 0 0 $X=322690 $Y=131520
X10317 1 2 DECAP5JI3V $T=329840 132160 1 180 $X=326610 $Y=131520
X10318 1 2 DECAP5JI3V $T=332080 42560 0 0 $X=331650 $Y=41920
X10319 1 2 DECAP5JI3V $T=333760 132160 0 0 $X=333330 $Y=131520
X10320 1 2 DECAP5JI3V $T=334320 105280 0 0 $X=333890 $Y=104640
X10321 1 2 DECAP5JI3V $T=352800 141120 1 180 $X=349570 $Y=140480
X10322 1 2 DECAP5JI3V $T=357840 132160 0 0 $X=357410 $Y=131520
X10323 1 2 DECAP5JI3V $T=357840 141120 1 0 $X=357410 $Y=136000
X10324 1 2 DECAP5JI3V $T=361200 42560 0 0 $X=360770 $Y=41920
X10325 1 2 DECAP5JI3V $T=361200 51520 1 0 $X=360770 $Y=46400
X10326 1 2 DECAP5JI3V $T=361200 159040 0 0 $X=360770 $Y=158400
X10327 1 2 DECAP5JI3V $T=366240 123200 0 0 $X=365810 $Y=122560
X10328 1 2 DECAP5JI3V $T=422240 24640 0 0 $X=421810 $Y=24000
X10329 1 2 DECAP5JI3V $T=422240 69440 1 0 $X=421810 $Y=64320
X10330 1 2 DECAP5JI3V $T=422240 78400 0 0 $X=421810 $Y=77760
X10331 1 2 DECAP5JI3V $T=422240 87360 0 0 $X=421810 $Y=86720
X10332 1 2 DECAP5JI3V $T=422240 96320 1 0 $X=421810 $Y=91200
X10333 1 2 DECAP5JI3V $T=422240 96320 0 0 $X=421810 $Y=95680
X10334 1 2 DECAP5JI3V $T=422240 105280 1 0 $X=421810 $Y=100160
X10335 1 2 DECAP5JI3V $T=422240 105280 0 0 $X=421810 $Y=104640
X10336 1 2 DECAP5JI3V $T=422240 114240 0 0 $X=421810 $Y=113600
X10337 1 2 DECAP5JI3V $T=422240 123200 1 0 $X=421810 $Y=118080
X10338 1 2 DECAP5JI3V $T=422240 132160 0 0 $X=421810 $Y=131520
X10339 1 2 DECAP5JI3V $T=422240 141120 1 0 $X=421810 $Y=136000
X10340 1 2 DECAP5JI3V $T=422240 150080 0 0 $X=421810 $Y=149440
X10341 1 2 DECAP5JI3V $T=422240 159040 1 0 $X=421810 $Y=153920
X10342 1 2 DECAP5JI3V $T=422240 176960 0 0 $X=421810 $Y=176320
X10343 1 2 DECAP5JI3V $T=422240 185920 1 0 $X=421810 $Y=180800
X10344 1 2 DECAP5JI3V $T=422240 194880 1 0 $X=421810 $Y=189760
X10345 1 2 DECAP5JI3V $T=422240 212800 0 0 $X=421810 $Y=212160
X10346 1 2 DECAP15JI3V $T=20160 33600 1 0 $X=19730 $Y=28480
X10347 1 2 DECAP15JI3V $T=20160 69440 0 0 $X=19730 $Y=68800
X10348 1 2 DECAP15JI3V $T=20160 123200 1 0 $X=19730 $Y=118080
X10349 1 2 DECAP15JI3V $T=20160 194880 1 0 $X=19730 $Y=189760
X10350 1 2 DECAP15JI3V $T=20160 203840 0 0 $X=19730 $Y=203200
X10351 1 2 DECAP15JI3V $T=34160 212800 0 0 $X=33730 $Y=212160
X10352 1 2 DECAP15JI3V $T=70000 33600 0 0 $X=69570 $Y=32960
X10353 1 2 DECAP15JI3V $T=75040 132160 0 0 $X=74610 $Y=131520
X10354 1 2 DECAP15JI3V $T=90720 123200 0 0 $X=90290 $Y=122560
X10355 1 2 DECAP15JI3V $T=100240 150080 0 0 $X=99810 $Y=149440
X10356 1 2 DECAP15JI3V $T=100240 159040 1 0 $X=99810 $Y=153920
X10357 1 2 DECAP15JI3V $T=100800 159040 0 0 $X=100370 $Y=158400
X10358 1 2 DECAP15JI3V $T=104720 114240 0 0 $X=104290 $Y=113600
X10359 1 2 DECAP15JI3V $T=104720 123200 1 0 $X=104290 $Y=118080
X10360 1 2 DECAP15JI3V $T=104720 185920 0 0 $X=104290 $Y=185280
X10361 1 2 DECAP15JI3V $T=104720 194880 1 0 $X=104290 $Y=189760
X10362 1 2 DECAP15JI3V $T=110320 212800 1 0 $X=109890 $Y=207680
X10363 1 2 DECAP15JI3V $T=110320 221760 1 0 $X=109890 $Y=216640
X10364 1 2 DECAP15JI3V $T=134400 87360 1 0 $X=133970 $Y=82240
X10365 1 2 DECAP15JI3V $T=134400 141120 1 0 $X=133970 $Y=136000
X10366 1 2 DECAP15JI3V $T=141120 78400 0 0 $X=140690 $Y=77760
X10367 1 2 DECAP15JI3V $T=148960 114240 1 0 $X=148530 $Y=109120
X10368 1 2 DECAP15JI3V $T=154000 221760 1 0 $X=153570 $Y=216640
X10369 1 2 DECAP15JI3V $T=177520 87360 1 0 $X=177090 $Y=82240
X10370 1 2 DECAP15JI3V $T=186480 78400 0 0 $X=186050 $Y=77760
X10371 1 2 DECAP15JI3V $T=206080 87360 0 0 $X=205650 $Y=86720
X10372 1 2 DECAP15JI3V $T=206080 150080 1 0 $X=205650 $Y=144960
X10373 1 2 DECAP15JI3V $T=206640 141120 1 0 $X=206210 $Y=136000
X10374 1 2 DECAP15JI3V $T=206640 159040 0 0 $X=206210 $Y=158400
X10375 1 2 DECAP15JI3V $T=206640 176960 0 0 $X=206210 $Y=176320
X10376 1 2 DECAP15JI3V $T=207760 96320 1 0 $X=207330 $Y=91200
X10377 1 2 DECAP15JI3V $T=208880 141120 0 0 $X=208450 $Y=140480
X10378 1 2 DECAP15JI3V $T=208880 203840 0 0 $X=208450 $Y=203200
X10379 1 2 DECAP15JI3V $T=210000 203840 1 0 $X=209570 $Y=198720
X10380 1 2 DECAP15JI3V $T=210560 221760 1 0 $X=210130 $Y=216640
X10381 1 2 DECAP15JI3V $T=211120 87360 1 0 $X=210690 $Y=82240
X10382 1 2 DECAP15JI3V $T=259280 96320 1 0 $X=258850 $Y=91200
X10383 1 2 DECAP15JI3V $T=270480 78400 0 0 $X=270050 $Y=77760
X10384 1 2 DECAP15JI3V $T=273840 114240 1 0 $X=273410 $Y=109120
X10385 1 2 DECAP15JI3V $T=279440 150080 0 0 $X=279010 $Y=149440
X10386 1 2 DECAP15JI3V $T=308560 123200 1 0 $X=308130 $Y=118080
X10387 1 2 DECAP15JI3V $T=308560 132160 1 0 $X=308130 $Y=127040
X10388 1 2 DECAP15JI3V $T=309680 87360 0 0 $X=309250 $Y=86720
X10389 1 2 DECAP15JI3V $T=309680 96320 1 0 $X=309250 $Y=91200
X10390 1 2 DECAP15JI3V $T=309680 123200 0 0 $X=309250 $Y=122560
X10391 1 2 DECAP15JI3V $T=311920 105280 0 0 $X=311490 $Y=104640
X10392 1 2 DECAP15JI3V $T=313600 114240 0 0 $X=313170 $Y=113600
X10393 1 2 DECAP15JI3V $T=316400 185920 1 0 $X=315970 $Y=180800
X10394 1 2 DECAP15JI3V $T=316960 51520 1 0 $X=316530 $Y=46400
X10395 1 2 DECAP15JI3V $T=316960 185920 0 0 $X=316530 $Y=185280
X10396 1 2 DECAP15JI3V $T=316960 194880 1 0 $X=316530 $Y=189760
X10397 1 2 DECAP15JI3V $T=332640 221760 1 0 $X=332210 $Y=216640
X10398 1 2 DECAP15JI3V $T=365120 176960 1 0 $X=364690 $Y=171840
X10399 1 2 DECAP15JI3V $T=366240 185920 0 0 $X=365810 $Y=185280
X10400 1 2 DECAP15JI3V $T=378560 78400 1 0 $X=378130 $Y=73280
X10401 1 2 DECAP15JI3V $T=379120 176960 1 0 $X=378690 $Y=171840
X10402 1 2 DECAP15JI3V $T=384720 42560 1 0 $X=384290 $Y=37440
X10403 1 2 DECAP15JI3V $T=384720 42560 0 0 $X=384290 $Y=41920
X10404 1 2 DECAP15JI3V $T=384720 168000 1 0 $X=384290 $Y=162880
X10405 1 2 DECAP15JI3V $T=400960 78400 1 0 $X=400530 $Y=73280
X10406 1 2 DECAP15JI3V $T=400960 87360 1 0 $X=400530 $Y=82240
X10407 1 2 DECAP15JI3V $T=400960 212800 1 0 $X=400530 $Y=207680
X10408 1 2 DECAP15JI3V $T=402080 185920 1 0 $X=401650 $Y=180800
X10409 1 2 DECAP15JI3V $T=404880 203840 0 0 $X=404450 $Y=203200
X10410 1 2 DECAP15JI3V $T=406000 176960 0 0 $X=405570 $Y=176320
X10411 1 2 DECAP15JI3V $T=408800 33600 1 0 $X=408370 $Y=28480
X10412 1 2 DECAP15JI3V $T=408800 114240 1 0 $X=408370 $Y=109120
X10413 1 2 DECAP15JI3V $T=408800 141120 0 0 $X=408370 $Y=140480
X10414 1 2 DECAP15JI3V $T=409920 96320 0 0 $X=409490 $Y=95680
X10415 1 2 DECAP15JI3V $T=409920 105280 1 0 $X=409490 $Y=100160
X10416 1 2 DECAP15JI3V $T=409920 114240 0 0 $X=409490 $Y=113600
X10417 1 2 DECAP15JI3V $T=409920 132160 0 0 $X=409490 $Y=131520
X10418 1 2 DECAP15JI3V $T=409920 141120 1 0 $X=409490 $Y=136000
X10419 1 2 DECAP15JI3V $T=416640 185920 0 0 $X=416210 $Y=185280
D0 83 1 p_ddnwmv AREA=8.4767e-08 PJ=0.00123324 perimeter=0.00123324 $X=17730 $Y=17520 $dt=2
D1 2 1 p_dipdnwmv AREA=1.66597e-09 PJ=0.000831805 perimeter=0.000831805 $X=27180 $Y=94080 $dt=3
D2 2 1 p_dipdnwmv AREA=1.65762e-09 PJ=0.000829452 perimeter=0.000829452 $X=28860 $Y=210560 $dt=3
D3 2 1 p_dipdnwmv AREA=1.66947e-09 PJ=0.000832178 perimeter=0.000832178 $X=40620 $Y=129920 $dt=3
D4 2 1 p_dipdnwmv AREA=1.65893e-09 PJ=0.000835699 perimeter=0.000835699 $X=53650 $Y=174710 $dt=3
D5 2 1 p_dipdnwmv AREA=1.6774e-09 PJ=0.000833895 perimeter=0.000833895 $X=57010 $Y=67190 $dt=3
D6 2 1 p_dipdnwmv AREA=1.62356e-09 PJ=0.000824013 perimeter=0.000824013 $X=91990 $Y=192430 $dt=3
D7 2 1 p_dipdnwmv AREA=1.66696e-09 PJ=0.000835085 perimeter=0.000835085 $X=101900 $Y=85110 $dt=3
D8 2 1 p_dipdnwmv AREA=1.65811e-09 PJ=0.000830245 perimeter=0.000830245 $X=101900 $Y=103030 $dt=3
D9 2 1 p_dipdnwmv AREA=1.66166e-09 PJ=0.000833269 perimeter=0.000833269 $X=101900 $Y=147830 $dt=3
D10 2 1 p_dipdnwmv AREA=1.6681e-09 PJ=0.000833335 perimeter=0.000833335 $X=113570 $Y=76150 $dt=3
D11 2 1 p_dipdnwmv AREA=1.66771e-09 PJ=0.000832586 perimeter=0.000832586 $X=118050 $Y=120950 $dt=3
D12 2 1 p_dipdnwmv AREA=1.6716e-09 PJ=0.000833709 perimeter=0.000833709 $X=143250 $Y=138870 $dt=3
D13 2 1 p_dipdnwmv AREA=1.66525e-09 PJ=0.000831652 perimeter=0.000831652 $X=143810 $Y=111990 $dt=3
D14 2 1 p_dipdnwmv AREA=1.67857e-09 PJ=0.000836374 perimeter=0.000836374 $X=144370 $Y=49270 $dt=3
D15 2 1 p_dipdnwmv AREA=1.67238e-09 PJ=0.000835208 perimeter=0.000835208 $X=146050 $Y=165750 $dt=3
D16 2 1 p_dipdnwmv AREA=1.66036e-09 PJ=0.000835202 perimeter=0.000835202 $X=161170 $Y=40310 $dt=3
D17 2 1 p_dipdnwmv AREA=1.67755e-09 PJ=0.000834786 perimeter=0.000834786 $X=164530 $Y=156790 $dt=3
D18 2 1 p_dipdnwmv AREA=1.08218e-09 PJ=0.000821773 perimeter=0.000821773 $X=164530 $Y=219510 $dt=3
D19 2 1 p_dipdnwmv AREA=1.6798e-09 PJ=0.000840932 perimeter=0.000840932 $X=179090 $Y=58230 $dt=3
D20 2 1 p_dipdnwmv AREA=1.6264e-09 PJ=0.000826294 perimeter=0.000826294 $X=189730 $Y=31350 $dt=3
D21 2 1 p_dipdnwmv AREA=1.6322e-09 PJ=0.00082472 perimeter=0.00082472 $X=207740 $Y=183670 $dt=3
D22 2 1 p_dipdnwmv AREA=1.61051e-09 PJ=0.000822069 perimeter=0.000822069 $X=273360 $Y=22480 $dt=3
D23 2 1 p_dipdnwmv AREA=1.63119e-09 PJ=0.000824905 perimeter=0.000824905 $X=273880 $Y=201390 $dt=3
.ends aska_dig

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: aska_dig_lvs                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt aska_dig_lvs gndd vdd3
** N=83 EP=2 FDC=26859
X0 vdd3 gndd 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70
+ 71 72 73 74 75 76 77 78 79 80
+ 81 82 aska_dig $T=9030 9935 0 0 $X=9110 $Y=9935
.ends aska_dig_lvs
