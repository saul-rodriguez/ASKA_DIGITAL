

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO aska_dig 
  PIN enable 
    ANTENNAPARTIALMETALAREA 0.3164 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.2769 LAYER MET3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA3 ;
    ANTENNADIFFAREA 1.6287 LAYER MET4 ; 
    ANTENNAPARTIALMETALAREA 61.4432 LAYER MET4 ;
    ANTENNAPARTIALMETALSIDEAREA 247.447 LAYER MET4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 7.89087 LAYER MET4 ; 
    ANTENNAMAXAREACAR 30.6269 LAYER MET4 ;
    ANTENNAMAXSIDEAREACAR 124.303 LAYER MET4 ;
    ANTENNAMAXCUTCAR 0.894994 LAYER VIATP ;
  END enable
  PIN pulse_active 
    ANTENNADIFFAREA 3.5375 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 2.5396 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.5655 LAYER MET3 ;
  END pulse_active
  PIN DAC[5] 
    ANTENNADIFFAREA 3.5375 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 1.396 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.6839 LAYER MET3 ;
  END DAC[5]
  PIN DAC[4] 
    ANTENNADIFFAREA 3.5375 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.304 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3334 LAYER MET3 ;
  END DAC[4]
  PIN DAC[3] 
    ANTENNADIFFAREA 3.5375 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.5236 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4295 LAYER MET3 ;
  END DAC[3]
  PIN DAC[2] 
    ANTENNADIFFAREA 3.5375 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.304 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3334 LAYER MET3 ;
  END DAC[2]
  PIN DAC[1] 
    ANTENNADIFFAREA 3.5375 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.252 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3334 LAYER MET3 ;
  END DAC[1]
  PIN DAC[0] 
    ANTENNADIFFAREA 3.5375 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.5236 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.4295 LAYER MET3 ;
  END DAC[0]
  PIN down_switches[31] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 46.4478 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 187.766 LAYER MET3 ;
  END down_switches[31]
  PIN down_switches[30] 
    ANTENNAPARTIALMETALAREA 0.9548 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8533 LAYER MET3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA3 ;
    ANTENNADIFFAREA 2.30485 LAYER MET4 ; 
    ANTENNAPARTIALMETALAREA 3.4808 LAYER MET4 ;
    ANTENNAPARTIALMETALSIDEAREA 13.9442 LAYER MET4 ;
  END down_switches[30]
  PIN down_switches[29] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 31.9788 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 129.057 LAYER MET3 ;
  END down_switches[29]
  PIN down_switches[28] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 37.7412 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 152.629 LAYER MET3 ;
  END down_switches[28]
  PIN down_switches[27] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 25.6788 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 103.949 LAYER MET3 ;
  END down_switches[27]
  PIN down_switches[26] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 25.1778 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 101.717 LAYER MET3 ;
  END down_switches[26]
  PIN down_switches[25] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 23.8 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 96.3664 LAYER MET3 ;
  END down_switches[25]
  PIN down_switches[24] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 15.7698 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 63.749 LAYER MET3 ;
  END down_switches[24]
  PIN down_switches[23] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.9548 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8533 LAYER MET3 ;
  END down_switches[23]
  PIN down_switches[22] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.3276 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3221 LAYER MET3 ;
  END down_switches[22]
  PIN down_switches[21] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 5.922 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.2159 LAYER MET3 ;
  END down_switches[21]
  PIN down_switches[20] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.1736 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7006 LAYER MET3 ;
  END down_switches[20]
  PIN down_switches[19] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.4844 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9549 LAYER MET3 ;
  END down_switches[19]
  PIN down_switches[18] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.4844 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9549 LAYER MET3 ;
  END down_switches[18]
  PIN down_switches[17] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.1736 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7006 LAYER MET3 ;
  END down_switches[17]
  PIN down_switches[16] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.4844 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9549 LAYER MET3 ;
  END down_switches[16]
  PIN down_switches[15] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.1736 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7006 LAYER MET3 ;
  END down_switches[15]
  PIN down_switches[14] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.4844 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9549 LAYER MET3 ;
  END down_switches[14]
  PIN down_switches[13] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.1402 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.35595 LAYER MET3 ;
  END down_switches[13]
  PIN down_switches[12] 
    ANTENNAPARTIALMETALAREA 0.6412 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.5877 LAYER MET3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA3 ;
    ANTENNADIFFAREA 2.30485 LAYER MET4 ; 
    ANTENNAPARTIALMETALAREA 2.2264 LAYER MET4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.8818 LAYER MET4 ;
  END down_switches[12]
  PIN down_switches[11] 
    ANTENNAPARTIALMETALAREA 0.1736 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7006 LAYER MET3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA3 ;
    ANTENNADIFFAREA 2.30485 LAYER MET4 ; 
    ANTENNAPARTIALMETALAREA 4.7352 LAYER MET4 ;
    ANTENNAPARTIALMETALSIDEAREA 19.0066 LAYER MET4 ;
  END down_switches[11]
  PIN down_switches[10] 
    ANTENNAPARTIALMETALAREA 0.9548 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8533 LAYER MET3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA3 ;
    ANTENNADIFFAREA 2.30485 LAYER MET4 ; 
    ANTENNAPARTIALMETALAREA 12.8888 LAYER MET4 ;
    ANTENNAPARTIALMETALSIDEAREA 51.9122 LAYER MET4 ;
  END down_switches[10]
  PIN down_switches[9] 
    ANTENNAPARTIALMETALAREA 0.9548 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8533 LAYER MET3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA3 ;
    ANTENNADIFFAREA 2.30485 LAYER MET4 ; 
    ANTENNAPARTIALMETALAREA 14.9272 LAYER MET4 ;
    ANTENNAPARTIALMETALSIDEAREA 60.1386 LAYER MET4 ;
  END down_switches[9]
  PIN down_switches[8] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 39.917 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 161.2 LAYER MET3 ;
  END down_switches[8]
  PIN down_switches[7] 
    ANTENNAPARTIALMETALAREA 0.1402 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.35595 LAYER MET3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA3 ;
    ANTENNADIFFAREA 2.30485 LAYER MET4 ; 
    ANTENNAPARTIALMETALAREA 2.9696 LAYER MET4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.091 LAYER MET4 ;
  END down_switches[7]
  PIN down_switches[6] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 42.3024 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 171.037 LAYER MET3 ;
  END down_switches[6]
  PIN down_switches[5] 
    ANTENNAPARTIALMETALAREA 0.1402 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.35595 LAYER MET3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA3 ;
    ANTENNADIFFAREA 2.30485 LAYER MET4 ; 
    ANTENNAPARTIALMETALAREA 1.7152 LAYER MET4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.0286 LAYER MET4 ;
  END down_switches[5]
  PIN down_switches[4] 
    ANTENNAPARTIALMETALAREA 0.1736 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7006 LAYER MET3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA3 ;
    ANTENNADIFFAREA 2.30485 LAYER MET4 ; 
    ANTENNAPARTIALMETALAREA 2.54 LAYER MET4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.1474 LAYER MET4 ;
  END down_switches[4]
  PIN down_switches[3] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 16.9148 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 68.2633 LAYER MET3 ;
  END down_switches[3]
  PIN down_switches[2] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 13.7508 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 55.8107 LAYER MET3 ;
  END down_switches[2]
  PIN down_switches[1] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 23.016 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 93.2024 LAYER MET3 ;
  END down_switches[1]
  PIN down_switches[0] 
    ANTENNADIFFAREA 2.30485 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 15.8004 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 64.0823 LAYER MET3 ;
  END down_switches[0]
  PIN up_switches[31] 
    ANTENNADIFFAREA 0.8862 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.3668 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7967 LAYER MET3 ;
  END up_switches[31]
  PIN up_switches[30] 
    ANTENNADIFFAREA 0.8862 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.304 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3334 LAYER MET3 ;
  END up_switches[30]
  PIN up_switches[29] 
    ANTENNADIFFAREA 0.8862 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.3668 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7967 LAYER MET3 ;
  END up_switches[29]
  PIN up_switches[28] 
    ANTENNADIFFAREA 0.8862 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.304 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3334 LAYER MET3 ;
  END up_switches[28]
  PIN up_switches[27] 
    ANTENNADIFFAREA 0.8862 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.3668 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7967 LAYER MET3 ;
  END up_switches[27]
  PIN up_switches[26] 
    ANTENNADIFFAREA 0.8862 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.6804 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0623 LAYER MET3 ;
  END up_switches[26]
  PIN up_switches[25] 
    ANTENNADIFFAREA 0.8862 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.6804 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0623 LAYER MET3 ;
  END up_switches[25]
  PIN up_switches[24] 
    ANTENNADIFFAREA 0.8862 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.8372 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6951 LAYER MET3 ;
  END up_switches[24]
  PIN up_switches[23] 
    ANTENNADIFFAREA 0.8862 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.3668 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7967 LAYER MET3 ;
  END up_switches[23]
  PIN up_switches[22] 
    ANTENNADIFFAREA 1.54144 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.1402 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.35595 LAYER MET3 ;
  END up_switches[22]
  PIN up_switches[21] 
    ANTENNADIFFAREA 0.8862 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.252 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3334 LAYER MET3 ;
  END up_switches[21]
  PIN up_switches[20] 
    ANTENNADIFFAREA 0.8862 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.3668 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7967 LAYER MET3 ;
  END up_switches[20]
  PIN up_switches[19] 
    ANTENNADIFFAREA 0.8862 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.304 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3334 LAYER MET3 ;
  END up_switches[19]
  PIN up_switches[18] 
    ANTENNADIFFAREA 1.6287 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.994 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3279 LAYER MET3 ;
  END up_switches[18]
  PIN up_switches[17] 
    ANTENNADIFFAREA 1.6287 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.994 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3279 LAYER MET3 ;
  END up_switches[17]
  PIN up_switches[16] 
    ANTENNADIFFAREA 1.6287 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 1.396 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.6839 LAYER MET3 ;
  END up_switches[16]
  PIN up_switches[15] 
    ANTENNADIFFAREA 1.6287 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.994 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3279 LAYER MET3 ;
  END up_switches[15]
  PIN up_switches[14] 
    ANTENNADIFFAREA 1.6287 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.994 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3279 LAYER MET3 ;
  END up_switches[14]
  PIN up_switches[13] 
    ANTENNADIFFAREA 1.6287 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.7212 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0171 LAYER MET3 ;
  END up_switches[13]
  PIN up_switches[12] 
    ANTENNADIFFAREA 1.6287 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 1.396 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.6839 LAYER MET3 ;
  END up_switches[12]
  PIN up_switches[11] 
    ANTENNADIFFAREA 1.6287 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 1.6016 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.78 LAYER MET3 ;
  END up_switches[11]
  PIN up_switches[10] 
    ANTENNADIFFAREA 1.6287 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.3668 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7967 LAYER MET3 ;
  END up_switches[10]
  PIN up_switches[9] 
    ANTENNADIFFAREA 1.6287 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.3668 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7967 LAYER MET3 ;
  END up_switches[9]
  PIN up_switches[8] 
    ANTENNADIFFAREA 1.6287 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.304 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3334 LAYER MET3 ;
  END up_switches[8]
  PIN up_switches[7] 
    ANTENNADIFFAREA 1.6287 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.252 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3334 LAYER MET3 ;
  END up_switches[7]
  PIN up_switches[6] 
    ANTENNADIFFAREA 1.6287 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.252 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3334 LAYER MET3 ;
  END up_switches[6]
  PIN up_switches[5] 
    ANTENNADIFFAREA 1.6287 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.8372 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6951 LAYER MET3 ;
  END up_switches[5]
  PIN up_switches[4] 
    ANTENNADIFFAREA 1.6287 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.6804 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.0623 LAYER MET3 ;
  END up_switches[4]
  PIN up_switches[3] 
    ANTENNADIFFAREA 1.54144 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.1736 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7006 LAYER MET3 ;
  END up_switches[3]
  PIN up_switches[2] 
    ANTENNADIFFAREA 1.54144 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.1736 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.7006 LAYER MET3 ;
  END up_switches[2]
  PIN up_switches[1] 
    ANTENNADIFFAREA 1.6287 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.304 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3334 LAYER MET3 ;
  END up_switches[1]
  PIN up_switches[0] 
    ANTENNADIFFAREA 1.6287 LAYER MET3 ; 
    ANTENNAPARTIALMETALAREA 0.304 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3334 LAYER MET3 ;
  END up_switches[0]
  PIN IC_addr[1] 
    ANTENNAPARTIALMETALAREA 0.4844 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9549 LAYER MET3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.954 LAYER MET3 ; 
    ANTENNAMAXAREACAR 9.14423 LAYER MET3 ;
    ANTENNAMAXSIDEAREACAR 37.3469 LAYER MET3 ;
    ANTENNAMAXCUTCAR 0.283438 LAYER VIA3 ;
  END IC_addr[1]
  PIN IC_addr[0] 
    ANTENNAPARTIALMETALAREA 3.5966 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.5149 LAYER MET3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.954 LAYER MET3 ; 
    ANTENNAMAXAREACAR 10.5927 LAYER MET3 ;
    ANTENNAMAXSIDEAREACAR 43.1923 LAYER MET3 ;
    ANTENNAMAXCUTCAR 0.283438 LAYER VIA3 ;
  END IC_addr[0]
  PIN SPI_MOSI 
    ANTENNAPARTIALMETALAREA 4.263 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.5206 LAYER MET3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.417 LAYER MET3 ; 
    ANTENNAMAXAREACAR 25.6638 LAYER MET3 ;
    ANTENNAMAXSIDEAREACAR 104.803 LAYER MET3 ;
    ANTENNAMAXCUTCAR 0.486331 LAYER VIA3 ;
  END SPI_MOSI
  PIN SPI_Clk 
    ANTENNAPARTIALMETALAREA 24.3528 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 98.2761 LAYER MET3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.417 LAYER MET3 ; 
    ANTENNAMAXAREACAR 60.66 LAYER MET3 ;
    ANTENNAMAXSIDEAREACAR 245.267 LAYER MET3 ;
    ANTENNAMAXCUTCAR 0.648441 LAYER VIA3 ;
  END SPI_Clk
  PIN SPI_CS 
    ANTENNAPARTIALMETALAREA 1.4762 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.96075 LAYER MET3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.774 LAYER MET3 ; 
    ANTENNAMAXAREACAR 18.7317 LAYER MET3 ;
    ANTENNAMAXSIDEAREACAR 76.6743 LAYER MET3 ;
    ANTENNAPARTIALCUTAREA 0.1352 LAYER VIA3 ;
    ANTENNAMAXCUTCAR 0.902742 LAYER VIA3 ;
    ANTENNAPARTIALMETALAREA 13.4752 LAYER MET4 ;
    ANTENNAPARTIALMETALSIDEAREA 54.4886 LAYER MET4 ;
    ANTENNAGATEAREA 17.835 LAYER MET4 ; 
    ANTENNAMAXAREACAR 19.4872 LAYER MET4 ;
    ANTENNAMAXSIDEAREACAR 79.7295 LAYER MET4 ;
    ANTENNAMAXCUTCAR 1.12528 LAYER VIATP ;
  END SPI_CS
  PIN porborn 
    ANTENNAPARTIALMETALAREA 0.994 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.3279 LAYER MET3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.417 LAYER MET3 ; 
    ANTENNAMAXAREACAR 19.0571 LAYER MET3 ;
    ANTENNAMAXSIDEAREACAR 77.6367 LAYER MET3 ;
    ANTENNAMAXCUTCAR 0.648441 LAYER VIA3 ;
  END porborn
  PIN reset_l 
    ANTENNAPARTIALMETALAREA 2.499 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.0853 LAYER MET3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6115 LAYER MET3 ; 
    ANTENNAMAXAREACAR 14.841 LAYER MET3 ;
    ANTENNAMAXSIDEAREACAR 60.2328 LAYER MET3 ;
    ANTENNAMAXCUTCAR 0.442191 LAYER VIA3 ;
  END reset_l
  PIN clk 
    ANTENNAPARTIALMETALAREA 23.1352 LAYER MET3 ;
    ANTENNAPARTIALMETALSIDEAREA 93.79 LAYER MET3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.54 LAYER MET3 ; 
    ANTENNAMAXAREACAR 44.4922 LAYER MET3 ;
    ANTENNAMAXSIDEAREACAR 180.706 LAYER MET3 ;
    ANTENNAMAXCUTCAR 0.500741 LAYER VIA3 ;
  END clk
END aska_dig

END LIBRARY
