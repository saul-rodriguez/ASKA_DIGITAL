* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : aska_dig                                     *
* Netlisted  : Mon Sep  9 14:22:33 2024                     *
* PVS Version: 23.10-p043 Mon Oct 2 18:09:08 PDT 2023      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(ne3i) nemi ndiff(D) p1trm(G) ndiff(S) pwitrm(B)
*.DEVTMPLT 1 MP(pe3i) pemi pdiff(D) p1trm(G) pdiff(S) dnwtrm(B)
*.DEVTMPLT 2 D(p_ddnwmv) p_ddnwmv bulk(POS) dnwtrm(NEG)
*.DEVTMPLT 3 D(p_dipdnwmv) p_dipwmv pwitrm(POS) dnwtrm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: EN2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt EN2JI3VX0 vdd3i! gnd3i! A B Q
*.DEVICECLIMB
** N=10 EP=5 FDC=10
M0 8 A 9 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=620 $Y=980 $dt=0
M1 gnd3i! B 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=1220 $Y=980 $dt=0
M2 7 A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=1.134e-13 PD=9.6e-07 PS=9.6e-07 $X=2110 $Y=980 $dt=0
M3 gnd3i! B 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.698e-13 AS=1.134e-13 PD=3.22e-06 PS=9.6e-07 $X=3000 $Y=980 $dt=0
M4 Q 9 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=2.058e-13 PD=1.8e-06 PS=1.82e-06 $X=4440 $Y=1020 $dt=0
M5 9 A vdd3i! vdd3i! pe3i L=3e-07 W=9e-07 AD=3.195e-13 AS=8.517e-13 PD=1.61e-06 PS=4.61e-06 $X=685 $Y=2410 $dt=1
M6 vdd3i! B 9 vdd3i! pe3i L=3e-07 W=9e-07 AD=4.30855e-13 AS=3.195e-13 PD=1.83273e-06 PS=1.61e-06 $X=1695 $Y=2410 $dt=1
M7 10 A vdd3i! vdd3i! pe3i L=3e-07 W=1.3e-06 AD=1.95e-13 AS=6.22345e-13 PD=1.6e-06 PS=2.64727e-06 $X=2825 $Y=2520 $dt=1
M8 Q B 10 vdd3i! pe3i L=3e-07 W=1.3e-06 AD=6.21324e-13 AS=1.95e-13 PD=2.52941e-06 PS=1.6e-06 $X=3425 $Y=2520 $dt=1
M9 vdd3i! 9 Q vdd3i! pe3i L=3e-07 W=9.1e-07 AD=8.0675e-13 AS=4.34926e-13 PD=4.39e-06 PS=1.77059e-06 $X=4575 $Y=2520 $dt=1
.ends EN2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO3JI3VX1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO3JI3VX1 vdd3i! gnd3i! C Q B A
*.DEVICECLIMB
** N=9 EP=6 FDC=6
M0 Q C gnd3i! gnd3i! ne3i L=3.4986e-07 W=8.92071e-07 AD=2.37813e-13 AS=4.30337e-13 PD=1.42707e-06 PS=2.76707e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! B Q gnd3i! ne3i L=3.4986e-07 W=8.92071e-07 AD=2.40287e-13 AS=2.37813e-13 PD=1.44207e-06 PS=1.42707e-06 $X=1500 $Y=660 $dt=0
M2 Q A gnd3i! gnd3i! ne3i L=3.4986e-07 W=8.92071e-07 AD=4.29162e-13 AS=2.40287e-13 PD=2.74707e-06 PS=1.44207e-06 $X=2390 $Y=660 $dt=0
M3 9 C vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=1.3994e-12 PD=1.72e-06 PS=5.15e-06 $X=955 $Y=2410 $dt=1
M4 8 B 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=2.1855e-13 PD=1.72e-06 PS=1.72e-06 $X=1565 $Y=2410 $dt=1
M5 Q A 8 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=2.1855e-13 PD=3.78e-06 PS=1.72e-06 $X=2175 $Y=2410 $dt=1
.ends NO3JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA2JI3VX2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA2JI3VX2 vdd3i! gnd3i! B Q A
*.DEVICECLIMB
** N=8 EP=5 FDC=8
M0 8 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=7.09e-13 PD=1.14e-06 PS=3.68e-06 $X=740 $Y=660 $dt=0
M1 Q A 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=1.1125e-13 PD=1.43e-06 PS=1.14e-06 $X=1340 $Y=660 $dt=0
M2 7 A Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=2.403e-13 PD=1.14e-06 PS=1.43e-06 $X=2230 $Y=660 $dt=0
M3 gnd3i! B 7 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=7.09e-13 AS=1.1125e-13 PD=3.68e-06 PS=1.14e-06 $X=2830 $Y=660 $dt=0
M4 Q B vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.7e-13 AS=8.172e-13 PD=1.54e-06 PS=4.22e-06 $X=540 $Y=2410 $dt=1
M5 vdd3i! A Q vdd3i! pe3i L=3e-07 W=1e-06 AD=8.172e-13 AS=2.7e-13 PD=4.22e-06 PS=1.54e-06 $X=1380 $Y=2410 $dt=1
M6 Q A vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.7e-13 AS=8.172e-13 PD=1.54e-06 PS=4.22e-06 $X=2240 $Y=2410 $dt=1
M7 vdd3i! B Q vdd3i! pe3i L=3e-07 W=1e-06 AD=8.172e-13 AS=2.7e-13 PD=4.22e-06 PS=1.54e-06 $X=3080 $Y=2410 $dt=1
.ends NA2JI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO22JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO22JI3VX1 vdd3i! gnd3i! B A Q C
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 8 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=4.87734e-13 PD=9.6e-07 PS=2.24324e-06 $X=720 $Y=1130 $dt=0
M1 gnd3i! A 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=4.87734e-13 AS=1.134e-13 PD=2.24324e-06 PS=9.6e-07 $X=1610 $Y=1130 $dt=0
M2 Q 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=1.03353e-12 PD=1.43e-06 PS=4.75353e-06 $X=2580 $Y=660 $dt=0
M3 gnd3i! C Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=6.098e-13 AS=2.403e-13 PD=3.52e-06 PS=1.43e-06 $X=3470 $Y=660 $dt=0
M4 10 B vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=1.0178e-12 PD=1.1e-06 PS=4.78e-06 $X=770 $Y=2410 $dt=1
M5 8 A 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.505e-13 AS=1.0625e-13 PD=2.76e-06 PS=1.1e-06 $X=1320 $Y=2410 $dt=1
M6 9 8 Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=6.768e-13 PD=1.66e-06 PS=3.78e-06 $X=2920 $Y=2410 $dt=1
M7 vdd3i! C 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=9.682e-13 AS=1.7625e-13 PD=4.66e-06 PS=1.66e-06 $X=3470 $Y=2410 $dt=1
.ends NO22JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DFRRQJI3VX2                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DFRRQJI3VX2 vdd3i! gnd3i! RN D C Q
*.DEVICECLIMB
** N=23 EP=6 FDC=32
M0 gnd3i! 17 19 gnd3i! ne3i L=3.5e-07 W=6.6e-07 AD=1.94849e-13 AS=3.168e-13 PD=1.21781e-06 PS=2.28e-06 $X=620 $Y=660 $dt=0
M1 10 RN gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.28952e-13 AS=2.62751e-13 PD=2.36956e-06 PS=1.64219e-06 $X=1510 $Y=660 $dt=0
M2 18 19 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.55236e-13 PD=6.7e-07 PS=1.11822e-06 $X=2340 $Y=1390 $dt=0
M3 17 9 18 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=2940 $Y=1390 $dt=0
M4 16 15 17 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=3830 $Y=1390 $dt=0
M5 10 D 16 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.835e-13 AS=5.25e-14 PD=2.19e-06 PS=6.7e-07 $X=4430 $Y=1390 $dt=0
M6 gnd3i! C 15 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.659e-13 AS=2.016e-13 PD=1.21e-06 PS=1.8e-06 $X=6060 $Y=1390 $dt=0
M7 9 15 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.95e-13 AS=1.659e-13 PD=2.23e-06 PS=1.21e-06 $X=7045 $Y=1390 $dt=0
M8 14 19 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=8695 $Y=1020 $dt=0
M9 13 9 14 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=9295 $Y=1020 $dt=0
M10 12 15 13 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=10185 $Y=1020 $dt=0
M11 8 11 12 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.55817e-13 AS=5.25e-14 PD=9.68244e-07 PS=6.7e-07 $X=10785 $Y=1020 $dt=0
M12 gnd3i! RN 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=5.94987e-13 AS=3.30183e-13 PD=3.35209e-06 PS=2.05176e-06 $X=11755 $Y=660 $dt=0
M13 11 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=6.6e-07 AD=3.168e-13 AS=4.41226e-13 PD=2.28e-06 PS=2.48582e-06 $X=12750 $Y=890 $dt=0
M14 Q 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=5.94987e-13 PD=1.43e-06 PS=3.35209e-06 $X=14380 $Y=660 $dt=0
M15 gnd3i! 13 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=2.403e-13 PD=2.74e-06 PS=1.43e-06 $X=15270 $Y=660 $dt=0
M16 vdd3i! 17 19 vdd3i! pe3i L=3e-07 W=1e-06 AD=2.97674e-13 AS=4.8e-13 PD=1.7907e-06 PS=2.96e-06 $X=620 $Y=2670 $dt=1
M17 17 RN vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.136e-13 AS=2.14326e-13 PD=2.4e-06 PS=1.2893e-06 $X=1460 $Y=2670 $dt=1
M18 23 19 vdd3i! vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=5.1875e-13 PD=6.7e-07 PS=2.99e-06 $X=3080 $Y=3400 $dt=1
M19 17 15 23 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=1.21617e-13 AS=5.25e-14 PD=9.13043e-07 PS=6.7e-07 $X=3630 $Y=3400 $dt=1
M20 22 9 17 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=1.2e-13 AS=2.77983e-13 PD=1.21e-06 PS=2.08696e-06 $X=4470 $Y=2860 $dt=1
M21 vdd3i! D 22 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=5.00229e-13 AS=1.2e-13 PD=2.34286e-06 PS=1.21e-06 $X=5020 $Y=2860 $dt=1
M22 15 C vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=4.56625e-13 AS=3.75171e-13 PD=2.86e-06 PS=1.75714e-06 $X=6060 $Y=2860 $dt=1
M23 vdd3i! 15 9 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.92547e-13 AS=3.528e-13 PD=1.8586e-06 PS=2.42e-06 $X=7720 $Y=2670 $dt=1
M24 21 19 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=1.25e-13 AS=5.45203e-13 PD=1.25e-06 PS=2.5814e-06 $X=8740 $Y=2820 $dt=1
M25 13 15 21 vdd3i! pe3i L=3e-07 W=1e-06 AD=2.96338e-13 AS=1.25e-13 PD=2.19718e-06 PS=1.25e-06 $X=9290 $Y=2820 $dt=1
M26 20 9 13 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=1.24462e-13 PD=6.7e-07 PS=9.22817e-07 $X=10150 $Y=3235 $dt=1
M27 vdd3i! 11 20 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=3.93439e-13 AS=5.25e-14 PD=1.64096e-06 PS=6.7e-07 $X=10700 $Y=3235 $dt=1
M28 vdd3i! RN 13 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=6.74468e-13 AS=2.976e-13 PD=2.81307e-06 PS=2.4e-06 $X=11900 $Y=2410 $dt=1
M29 11 13 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=4.8e-13 AS=9.36761e-13 PD=2.96e-06 PS=3.90704e-06 $X=12740 $Y=2410 $dt=1
M30 Q 13 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=1.32083e-12 PD=1.95e-06 PS=5.50893e-06 $X=14440 $Y=2410 $dt=1
M31 vdd3i! 13 Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=8.802e-13 AS=3.807e-13 PD=4.56e-06 PS=1.95e-06 $X=15280 $Y=2410 $dt=1
.ends DFRRQJI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX8                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX8 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=19
M0 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=6.098e-13 PD=1.43e-06 PS=3.52e-06 $X=660 $Y=660 $dt=0
M1 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.804e-13 AS=2.403e-13 PD=1.91e-06 PS=1.43e-06 $X=1550 $Y=660 $dt=0
M2 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.804e-13 PD=1.43e-06 PS=1.91e-06 $X=2570 $Y=660 $dt=0
M3 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=3460 $Y=660 $dt=0
M4 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=4430 $Y=660 $dt=0
M5 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=5320 $Y=660 $dt=0
M6 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=6290 $Y=660 $dt=0
M7 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=8.702e-13 AS=2.403e-13 PD=3.94e-06 PS=1.43e-06 $X=7180 $Y=660 $dt=0
M8 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=5.51013e-13 PD=1.86506e-06 PS=3.69506e-06 $X=620 $Y=2410 $dt=1
M9 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.61963e-13 AS=2.83187e-13 PD=1.87506e-06 PS=1.86506e-06 $X=1170 $Y=2410 $dt=1
M10 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.61963e-13 PD=1.86506e-06 PS=1.87506e-06 $X=2020 $Y=2410 $dt=1
M11 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.61963e-13 AS=2.83187e-13 PD=1.87506e-06 PS=1.86506e-06 $X=2570 $Y=2410 $dt=1
M12 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.61963e-13 PD=1.86506e-06 PS=1.87506e-06 $X=3420 $Y=2410 $dt=1
M13 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.61963e-13 AS=2.83187e-13 PD=1.87506e-06 PS=1.86506e-06 $X=3970 $Y=2410 $dt=1
M14 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.61963e-13 PD=1.86506e-06 PS=1.87506e-06 $X=4820 $Y=2410 $dt=1
M15 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.61963e-13 AS=2.83187e-13 PD=1.87506e-06 PS=1.86506e-06 $X=5370 $Y=2410 $dt=1
M16 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.61963e-13 PD=1.86506e-06 PS=1.87506e-06 $X=6220 $Y=2410 $dt=1
M17 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.61963e-13 AS=2.83187e-13 PD=1.87506e-06 PS=1.86506e-06 $X=6770 $Y=2410 $dt=1
M18 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=5.79287e-13 AS=2.61963e-13 PD=3.69506e-06 PS=1.87506e-06 $X=7620 $Y=2410 $dt=1
.ends BUJI3VX8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DFRRQJI3VX4                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DFRRQJI3VX4 vdd3i! gnd3i! RN D C Q
*.DEVICECLIMB
** N=23 EP=6 FDC=36
M0 gnd3i! 17 19 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=4.272e-13 PD=1.43e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 10 RN gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.28952e-13 AS=2.403e-13 PD=2.36956e-06 PS=1.43e-06 $X=1510 $Y=660 $dt=0
M2 18 19 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.55236e-13 PD=6.7e-07 PS=1.11822e-06 $X=2340 $Y=1390 $dt=0
M3 17 9 18 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=2940 $Y=1390 $dt=0
M4 16 15 17 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=3830 $Y=1390 $dt=0
M5 10 D 16 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.835e-13 AS=5.25e-14 PD=2.19e-06 PS=6.7e-07 $X=4430 $Y=1390 $dt=0
M6 gnd3i! C 15 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.659e-13 AS=2.016e-13 PD=1.21e-06 PS=1.8e-06 $X=6060 $Y=1390 $dt=0
M7 9 15 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.95e-13 AS=1.659e-13 PD=2.23e-06 PS=1.21e-06 $X=7045 $Y=1390 $dt=0
M8 14 19 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=8695 $Y=1020 $dt=0
M9 13 9 14 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=9295 $Y=1020 $dt=0
M10 12 15 13 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=10185 $Y=1020 $dt=0
M11 8 11 12 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.55817e-13 AS=5.25e-14 PD=9.68244e-07 PS=6.7e-07 $X=10785 $Y=1020 $dt=0
M12 gnd3i! RN 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.60325e-13 AS=3.30183e-13 PD=1.475e-06 PS=2.05176e-06 $X=11755 $Y=660 $dt=0
M13 11 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=2.60325e-13 PD=2.74e-06 PS=1.475e-06 $X=12690 $Y=660 $dt=0
M14 Q 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=4.272e-13 PD=1.43e-06 PS=2.74e-06 $X=14280 $Y=660 $dt=0
M15 gnd3i! 13 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=15170 $Y=660 $dt=0
M16 Q 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=16060 $Y=660 $dt=0
M17 gnd3i! 13 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=2.403e-13 PD=2.74e-06 PS=1.43e-06 $X=16950 $Y=660 $dt=0
M18 vdd3i! 17 19 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.54046e-13 AS=6.768e-13 PD=2.58169e-06 PS=3.78e-06 $X=620 $Y=2410 $dt=1
M19 17 RN vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.136e-13 AS=2.31854e-13 PD=2.4e-06 PS=1.31831e-06 $X=1460 $Y=2670 $dt=1
M20 23 19 vdd3i! vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=5.1875e-13 PD=6.7e-07 PS=2.99e-06 $X=3080 $Y=3400 $dt=1
M21 17 15 23 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=1.21617e-13 AS=5.25e-14 PD=9.13043e-07 PS=6.7e-07 $X=3630 $Y=3400 $dt=1
M22 22 9 17 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=1.2e-13 AS=2.77983e-13 PD=1.21e-06 PS=2.08696e-06 $X=4470 $Y=2860 $dt=1
M23 vdd3i! D 22 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=5.00229e-13 AS=1.2e-13 PD=2.34286e-06 PS=1.21e-06 $X=5020 $Y=2860 $dt=1
M24 15 C vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=4.94875e-13 AS=3.75171e-13 PD=3.04e-06 PS=1.75714e-06 $X=6060 $Y=2860 $dt=1
M25 vdd3i! 15 9 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.92547e-13 AS=3.528e-13 PD=1.8586e-06 PS=2.42e-06 $X=7720 $Y=2670 $dt=1
M26 21 19 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=1.25e-13 AS=5.45203e-13 PD=1.25e-06 PS=2.5814e-06 $X=8740 $Y=2820 $dt=1
M27 13 15 21 vdd3i! pe3i L=3e-07 W=1e-06 AD=2.96338e-13 AS=1.25e-13 PD=2.19718e-06 PS=1.25e-06 $X=9290 $Y=2820 $dt=1
M28 20 9 13 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=1.24462e-13 PD=6.7e-07 PS=9.22817e-07 $X=10150 $Y=3235 $dt=1
M29 vdd3i! 11 20 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=2.90656e-13 AS=5.25e-14 PD=1.25671e-06 PS=6.7e-07 $X=10700 $Y=3235 $dt=1
M30 vdd3i! RN 13 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=4.98268e-13 AS=2.976e-13 PD=2.15435e-06 PS=2.4e-06 $X=11900 $Y=2410 $dt=1
M31 11 13 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=9.75775e-13 PD=3.78e-06 PS=4.21894e-06 $X=12740 $Y=2410 $dt=1
M32 Q 13 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=1.1618e-12 PD=1.95e-06 PS=4.88e-06 $X=14480 $Y=2410 $dt=1
M33 vdd3i! 13 Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=3.807e-13 PD=1.95e-06 PS=1.95e-06 $X=15320 $Y=2410 $dt=1
M34 Q 13 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=3.807e-13 PD=1.95e-06 PS=1.95e-06 $X=16160 $Y=2410 $dt=1
M35 vdd3i! 13 Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=3.807e-13 PD=3.78e-06 PS=1.95e-06 $X=17000 $Y=2410 $dt=1
.ends DFRRQJI3VX4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX1 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=4
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.44533e-13 AS=2.016e-13 PD=1.44667e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=6.6e-07 AD=2.88e-13 AS=3.84267e-13 PD=2.28e-06 PS=2.27333e-06 $X=1590 $Y=890 $dt=0
M2 vdd3i! A 6 vdd3i! pe3i L=3e-07 W=9e-07 AD=4.7931e-13 AS=4.32e-13 PD=1.95649e-06 PS=2.76e-06 $X=620 $Y=2410 $dt=1
M3 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=5.712e-13 AS=7.7739e-13 PD=3.70971e-06 PS=3.17322e-06 $X=1640 $Y=2410 $dt=1
.ends BUJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO3I2JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO3I2JI3VX1 vdd3i! gnd3i! AN BN C Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 8 AN 9 gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=6e-14 AS=2.304e-13 PD=7.3e-07 PS=1.92e-06 $X=620 $Y=1070 $dt=0
M1 gnd3i! BN 8 gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=1.98937e-13 AS=6e-14 PD=1.31617e-06 PS=7.3e-07 $X=1220 $Y=1070 $dt=0
M2 Q C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.68863e-13 PD=1.43e-06 PS=2.4404e-06 $X=2060 $Y=660 $dt=0
M3 gnd3i! 9 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.329e-13 AS=2.403e-13 PD=2.77e-06 PS=1.43e-06 $X=2950 $Y=660 $dt=0
M4 9 AN vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=5.71409e-13 PD=1.24e-06 PS=2.5758e-06 $X=560 $Y=2590 $dt=1
M5 vdd3i! BN 9 vdd3i! pe3i L=3e-07 W=7e-07 AD=5.71409e-13 AS=1.89e-13 PD=2.5758e-06 PS=1.24e-06 $X=1400 $Y=2590 $dt=1
M6 10 C vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=1.15098e-12 PD=1.66e-06 PS=5.1884e-06 $X=2330 $Y=2410 $dt=1
M7 Q 9 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=8.46e-13 AS=1.7625e-13 PD=4.02e-06 PS=1.66e-06 $X=2880 $Y=2410 $dt=1
.ends NO3I2JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: FAJI3VX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt FAJI3VX1 vdd3i! gnd3i! S CI B A CO
*.DEVICECLIMB
** N=20 EP=7 FDC=28
M0 gnd3i! 12 S gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.361e-13 AS=4.272e-13 PD=2.76e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 15 CI 12 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=7.375e-14 AS=2.832e-13 PD=8.4e-07 PS=2.14e-06 $X=2220 $Y=960 $dt=0
M2 14 B 15 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=7.375e-14 AS=7.375e-14 PD=8.4e-07 PS=8.4e-07 $X=2820 $Y=960 $dt=0
M3 gnd3i! A 14 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=2.34033e-13 AS=7.375e-14 PD=1.52158e-06 PS=8.4e-07 $X=3420 $Y=960 $dt=0
M4 13 CI gnd3i! gnd3i! ne3i L=3.5e-07 W=5.5e-07 AD=1.485e-13 AS=2.18167e-13 PD=1.09e-06 PS=1.41842e-06 $X=4350 $Y=660 $dt=0
M5 gnd3i! A 13 gnd3i! ne3i L=3.5e-07 W=5.5e-07 AD=2.5017e-13 AS=1.485e-13 PD=1.58058e-06 PS=1.09e-06 $X=5240 $Y=660 $dt=0
M6 13 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=1.296e-13 AS=2.1833e-13 PD=1.02e-06 PS=1.37942e-06 $X=6220 $Y=960 $dt=0
M7 12 10 13 gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=2.304e-13 AS=1.296e-13 PD=1.92e-06 PS=1.02e-06 $X=7110 $Y=960 $dt=0
M8 gnd3i! 10 CO gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=3.345e-13 AS=2.832e-13 PD=1.73e-06 PS=2.14e-06 $X=8700 $Y=960 $dt=0
M9 11 A gnd3i! gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=7.375e-14 AS=3.345e-13 PD=8.4e-07 PS=1.73e-06 $X=9830 $Y=960 $dt=0
M10 10 B 11 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=1.593e-13 AS=7.375e-14 PD=1.13e-06 PS=8.4e-07 $X=10430 $Y=960 $dt=0
M11 9 CI 10 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=1.593e-13 AS=1.593e-13 PD=1.13e-06 PS=1.13e-06 $X=11320 $Y=960 $dt=0
M12 gnd3i! B 9 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=4.382e-13 AS=1.593e-13 PD=1.95e-06 PS=1.13e-06 $X=12210 $Y=960 $dt=0
M13 9 A gnd3i! gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=3.068e-13 AS=4.382e-13 PD=2.22e-06 PS=1.95e-06 $X=13550 $Y=960 $dt=0
M14 vdd3i! 12 S vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.6395e-13 AS=7.1205e-13 PD=4.52213e-06 PS=3.83e-06 $X=645 $Y=2410 $dt=1
M15 vdd3i! CI 17 vdd3i! pe3i L=3e-07 W=1.03e-06 AD=4.8155e-13 AS=4.79437e-13 PD=2.35e-06 PS=3.03778e-06 $X=2125 $Y=2490 $dt=1
M16 17 B vdd3i! vdd3i! pe3i L=3e-07 W=1.03e-06 AD=3.0385e-13 AS=4.8155e-13 PD=1.62e-06 PS=2.35e-06 $X=3095 $Y=2490 $dt=1
M17 vdd3i! A 17 vdd3i! pe3i L=3e-07 W=1.03e-06 AD=4.1015e-13 AS=3.0385e-13 PD=2.01e-06 PS=1.62e-06 $X=3985 $Y=2490 $dt=1
M18 20 A vdd3i! vdd3i! pe3i L=3e-07 W=1.03e-06 AD=1.545e-13 AS=4.1015e-13 PD=1.33e-06 PS=2.01e-06 $X=4955 $Y=2490 $dt=1
M19 19 B 20 vdd3i! pe3i L=3e-07 W=1.03e-06 AD=1.545e-13 AS=1.545e-13 PD=1.33e-06 PS=1.33e-06 $X=5555 $Y=2490 $dt=1
M20 12 CI 19 vdd3i! pe3i L=3e-07 W=1.03e-06 AD=3.0385e-13 AS=1.545e-13 PD=1.62e-06 PS=1.33e-06 $X=6155 $Y=2490 $dt=1
M21 17 10 12 vdd3i! pe3i L=3e-07 W=1.03e-06 AD=6.9155e-13 AS=3.0385e-13 PD=3.77e-06 PS=1.62e-06 $X=7045 $Y=2490 $dt=1
M22 vdd3i! 10 CO vdd3i! pe3i L=3e-07 W=1.11e-06 AD=4.54624e-13 AS=5.6055e-13 PD=2.27286e-06 PS=3.23e-06 $X=8675 $Y=2410 $dt=1
M23 16 A vdd3i! vdd3i! pe3i L=3e-07 W=9.9e-07 AD=2.9205e-13 AS=4.05476e-13 PD=1.58e-06 PS=2.02714e-06 $X=9645 $Y=2530 $dt=1
M24 vdd3i! B 16 vdd3i! pe3i L=3e-07 W=9.9e-07 AD=5.763e-13 AS=2.9205e-13 PD=3.59e-06 PS=1.58e-06 $X=10535 $Y=2530 $dt=1
M25 10 CI 16 vdd3i! pe3i L=3e-07 W=1e-06 AD=2.95e-13 AS=4.65e-13 PD=1.59e-06 PS=3.01e-06 $X=12085 $Y=2520 $dt=1
M26 18 B 10 vdd3i! pe3i L=3e-07 W=1e-06 AD=1.5e-13 AS=2.95e-13 PD=1.3e-06 PS=1.59e-06 $X=12975 $Y=2520 $dt=1
M27 vdd3i! A 18 vdd3i! pe3i L=3e-07 W=1e-06 AD=8.18e-13 AS=1.5e-13 PD=4.39e-06 PS=1.3e-06 $X=13575 $Y=2520 $dt=1
.ends FAJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OR2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OR2JI3VX0 vdd3i! gnd3i! A B Q
*.DEVICECLIMB
** N=8 EP=5 FDC=6
M0 7 A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.75467e-13 PD=9.6e-07 PS=2.95333e-06 $X=530 $Y=1130 $dt=0
M1 gnd3i! B 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.75467e-13 AS=1.134e-13 PD=2.95333e-06 PS=9.6e-07 $X=1420 $Y=1130 $dt=0
M2 Q 7 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=5.75467e-13 PD=1.8e-06 PS=2.95333e-06 $X=2390 $Y=1130 $dt=0
M3 8 A 7 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=4.08e-13 PD=1.1e-06 PS=2.66e-06 $X=620 $Y=2410 $dt=1
M4 vdd3i! B 8 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=8.28174e-13 AS=1.0625e-13 PD=2.99419e-06 PS=1.1e-06 $X=1170 $Y=2410 $dt=1
M5 Q 7 vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=3.36e-13 AS=6.82026e-13 PD=2.36e-06 PS=2.46581e-06 $X=2440 $Y=2410 $dt=1
.ends OR2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA3I1JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA3I1JI3VX1 vdd3i! gnd3i! AN Q B C
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 gnd3i! AN 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.40779e-13 AS=2.016e-13 PD=1.24397e-06 PS=1.8e-06 $X=620 $Y=660 $dt=0
M1 9 10 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.26825e-13 AS=5.10221e-13 PD=1.175e-06 PS=2.63603e-06 $X=1670 $Y=660 $dt=0
M2 8 B 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.31275e-13 AS=1.26825e-13 PD=1.185e-06 PS=1.175e-06 $X=2305 $Y=660 $dt=0
M3 Q C 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=1.31275e-13 PD=2.74e-06 PS=1.185e-06 $X=2950 $Y=660 $dt=0
M4 vdd3i! AN 10 vdd3i! pe3i L=3e-07 W=7e-07 AD=4.82246e-13 AS=3.36e-13 PD=2.26063e-06 PS=2.36e-06 $X=620 $Y=2410 $dt=1
M5 vdd3i! 10 Q vdd3i! pe3i L=3.00059e-07 W=1.00314e-06 AD=6.91085e-13 AS=2.195e-13 PD=3.2396e-06 PS=1.46314e-06 $X=1430 $Y=2410 $dt=1
M6 Q B vdd3i! vdd3i! pe3i L=3.00059e-07 W=1.00314e-06 AD=2.195e-13 AS=6.91085e-13 PD=1.46314e-06 PS=3.2396e-06 $X=2270 $Y=2410 $dt=1
M7 Q C vdd3i! vdd3i! pe3i L=3.00059e-07 W=1.00314e-06 AD=4.232e-13 AS=6.91085e-13 PD=2.85314e-06 PS=3.2396e-06 $X=3000 $Y=2410 $dt=1
.ends NA3I1JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DLY2JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DLY2JI3VX1 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=12 EP=4 FDC=12
M0 gnd3i! A 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.577e-13 AS=2.016e-13 PD=1.79e-06 PS=1.8e-06 $X=620 $Y=660 $dt=0
M1 8 10 gnd3i! gnd3i! ne3i L=8e-07 W=4.2e-07 AD=2.548e-13 AS=3.577e-13 PD=1.7e-06 PS=1.79e-06 $X=1990 $Y=660 $dt=0
M2 8 10 9 gnd3i! ne3i L=8e-07 W=4.2e-07 AD=2.548e-13 AS=2.016e-13 PD=1.7e-06 PS=1.8e-06 $X=1990 $Y=1360 $dt=0
M3 gnd3i! 9 7 gnd3i! ne3i L=1e-06 W=4.2e-07 AD=3.42444e-13 AS=2.1e-13 PD=1.66718e-06 PS=1.62e-06 $X=3950 $Y=660 $dt=0
M4 6 9 7 gnd3i! ne3i L=1e-06 W=4.2e-07 AD=2.10588e-13 AS=2.1e-13 PD=1.81778e-06 PS=1.62e-06 $X=3950 $Y=1360 $dt=0
M5 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=7.25656e-13 PD=2.74e-06 PS=3.53282e-06 $X=6310 $Y=660 $dt=0
M6 vdd3i! A 10 vdd3i! pe3i L=3e-07 W=7e-07 AD=5.42937e-13 AS=3.535e-13 PD=2.69375e-06 PS=2.41e-06 $X=645 $Y=3120 $dt=1
M7 12 10 9 vdd3i! pe3i L=7.4e-07 W=4.2e-07 AD=2.8095e-13 AS=2.0035e-13 PD=1.785e-06 PS=1.77071e-06 $X=2050 $Y=2640 $dt=1
M8 12 10 vdd3i! vdd3i! pe3i L=7.4e-07 W=4.2e-07 AD=2.8095e-13 AS=3.25762e-13 PD=1.785e-06 PS=1.61625e-06 $X=2050 $Y=3400 $dt=1
M9 6 9 11 vdd3i! pe3i L=1e-06 W=4.2e-07 AD=2.856e-13 AS=2.479e-13 PD=2.2e-06 PS=1.715e-06 $X=4030 $Y=2660 $dt=1
M10 vdd3i! 9 11 vdd3i! pe3i L=1e-06 W=4.2e-07 AD=2.62018e-13 AS=2.479e-13 PD=1.40689e-06 PS=1.715e-06 $X=4030 $Y=3400 $dt=1
M11 Q 6 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.1205e-13 AS=8.79632e-13 PD=3.83e-06 PS=4.72311e-06 $X=6335 $Y=2410 $dt=1
.ends DLY2JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA3JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA3JI3VX0 vdd3i! gnd3i! C Q B A
*.DEVICECLIMB
** N=9 EP=6 FDC=6
M0 9 C gnd3i! gnd3i! ne3i L=3.5e-07 W=7e-07 AD=8.75e-14 AS=5.605e-13 PD=9.5e-07 PS=3.52e-06 $X=630 $Y=850 $dt=0
M1 8 B 9 gnd3i! ne3i L=3.5e-07 W=7e-07 AD=8.75e-14 AS=8.75e-14 PD=9.5e-07 PS=9.5e-07 $X=1230 $Y=850 $dt=0
M2 Q A 8 gnd3i! ne3i L=3.5e-07 W=7e-07 AD=3.36e-13 AS=8.75e-14 PD=2.36e-06 PS=9.5e-07 $X=1830 $Y=850 $dt=0
M3 Q C vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=5.76467e-13 PD=1.24e-06 PS=3.21333e-06 $X=470 $Y=2580 $dt=1
M4 vdd3i! B Q vdd3i! pe3i L=3e-07 W=7e-07 AD=5.76467e-13 AS=1.89e-13 PD=3.21333e-06 PS=1.24e-06 $X=1310 $Y=2580 $dt=1
M5 Q A vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=4.708e-13 AS=5.76467e-13 PD=3.92e-06 PS=3.21333e-06 $X=2040 $Y=2470 $dt=1
.ends NA3JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ON21JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ON21JI3VX1 vdd3i! gnd3i! B A Q C
*.DEVICECLIMB
** N=9 EP=6 FDC=6
M0 gnd3i! B 8 gnd3i! ne3i L=3.4958e-07 W=8.92071e-07 AD=2.40125e-13 AS=4.24712e-13 PD=1.43207e-06 PS=2.73707e-06 $X=615 $Y=660 $dt=0
M1 8 A gnd3i! gnd3i! ne3i L=3.4958e-07 W=8.92071e-07 AD=2.37987e-13 AS=2.40125e-13 PD=1.42707e-06 PS=1.43207e-06 $X=1505 $Y=660 $dt=0
M2 Q C 8 gnd3i! ne3i L=3.4958e-07 W=8.92071e-07 AD=4.24712e-13 AS=2.37987e-13 PD=2.73707e-06 PS=1.42707e-06 $X=2395 $Y=660 $dt=0
M3 9 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=9.418e-13 PD=1.66e-06 PS=4.63e-06 $X=695 $Y=2410 $dt=1
M4 Q A 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.75706e-13 AS=1.7625e-13 PD=2.44322e-06 PS=1.66e-06 $X=1245 $Y=2410 $dt=1
M5 vdd3i! C Q vdd3i! pe3i L=3e-07 W=9.85e-07 AD=1.1721e-12 AS=3.32319e-13 PD=4.94e-06 PS=1.70678e-06 $X=2210 $Y=2410 $dt=1
.ends ON21JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OA21JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OA21JI3VX1 vdd3i! gnd3i! C A B Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 8 C 9 gnd3i! ne3i L=3.5e-07 W=5.4e-07 AD=3.313e-13 AS=2.97e-13 PD=1.95333e-06 PS=2.18e-06 $X=690 $Y=660 $dt=0
M1 8 A gnd3i! gnd3i! ne3i L=3.5e-07 W=5.4e-07 AD=3.313e-13 AS=2.592e-13 PD=1.95333e-06 PS=2.04e-06 $X=1620 $Y=1480 $dt=0
M2 gnd3i! B 8 gnd3i! ne3i L=3.5e-07 W=5.4e-07 AD=2.92808e-13 AS=3.313e-13 PD=1.47273e-06 PS=1.95333e-06 $X=2450 $Y=1010 $dt=0
M3 Q 9 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=4.82592e-13 PD=2.74e-06 PS=2.42727e-06 $X=3510 $Y=660 $dt=0
M4 9 C vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=2.295e-13 AS=1.03315e-12 PD=1.39e-06 PS=4.25e-06 $X=975 $Y=2880 $dt=1
M5 10 A 9 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=2.295e-13 PD=1.1e-06 PS=1.39e-06 $X=1815 $Y=2880 $dt=1
M6 vdd3i! B 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.77448e-13 AS=1.0625e-13 PD=1.94425e-06 PS=1.1e-06 $X=2365 $Y=2880 $dt=1
M7 Q 9 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=7.92002e-13 PD=3.78e-06 PS=3.22516e-06 $X=3560 $Y=2410 $dt=1
.ends OA21JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX3                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX3 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=7
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=5.23e-13 AS=4.272e-13 PD=2.14e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.5365e-13 AS=5.23e-13 PD=1.46e-06 PS=2.14e-06 $X=1870 $Y=660 $dt=0
M2 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=7.586e-13 AS=2.5365e-13 PD=3.76e-06 PS=1.46e-06 $X=2790 $Y=660 $dt=0
M3 vdd3i! A 6 vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=6.11825e-13 AS=5.712e-13 PD=2.51971e-06 PS=3.70971e-06 $X=620 $Y=2410 $dt=1
M4 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=6.11825e-13 PD=1.87971e-06 PS=2.51971e-06 $X=1510 $Y=2410 $dt=1
M5 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=3.3675e-13 AS=2.751e-13 PD=1.92971e-06 PS=1.87971e-06 $X=2350 $Y=2410 $dt=1
M6 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=5.712e-13 AS=3.3675e-13 PD=3.70971e-06 PS=1.92971e-06 $X=3000 $Y=2410 $dt=1
.ends BUJI3VX3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AN211JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AN211JI3VX1 vdd3i! gnd3i! B A Q C D
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 9 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=6.47e-13 PD=1.14e-06 PS=3.58e-06 $X=690 $Y=660 $dt=0
M1 Q A 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.9785e-13 AS=1.1125e-13 PD=1.71704e-06 PS=1.14e-06 $X=1290 $Y=660 $dt=0
M2 gnd3i! C Q gnd3i! ne3i L=3.5e-07 W=6.65e-07 AD=5.036e-13 AS=2.2255e-13 PD=2.145e-06 PS=1.28296e-06 $X=2250 $Y=885 $dt=0
M3 Q D gnd3i! gnd3i! ne3i L=3.5e-07 W=6.65e-07 AD=3.22525e-13 AS=5.036e-13 PD=2.3e-06 PS=2.145e-06 $X=3505 $Y=885 $dt=0
M4 vdd3i! B 11 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.5825e-13 AS=6.768e-13 PD=2.06e-06 PS=3.78e-06 $X=620 $Y=2410 $dt=1
M5 11 A vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=4.5825e-13 PD=2e-06 PS=2.06e-06 $X=1570 $Y=2410 $dt=1
M6 10 C 11 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.115e-13 AS=4.1595e-13 PD=1.71e-06 PS=2e-06 $X=2460 $Y=2410 $dt=1
M7 Q D 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=2.115e-13 PD=3.78e-06 PS=1.71e-06 $X=3060 $Y=2410 $dt=1
.ends AN211JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX16                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX16 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=39
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=4.272e-13 PD=1.43e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=1510 $Y=660 $dt=0
M2 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=2400 $Y=660 $dt=0
M3 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=3290 $Y=660 $dt=0
M4 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=4180 $Y=660 $dt=0
M5 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.4475e-13 AS=2.403e-13 PD=1.44e-06 PS=1.43e-06 $X=5070 $Y=660 $dt=0
M6 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.63267e-13 AS=2.4475e-13 PD=1.95905e-06 PS=1.44e-06 $X=5970 $Y=660 $dt=0
M7 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.26533e-13 PD=1.34e-06 PS=1.76095e-06 $X=6940 $Y=750 $dt=0
M8 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=7830 $Y=750 $dt=0
M9 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=8800 $Y=750 $dt=0
M10 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=9690 $Y=750 $dt=0
M11 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=10660 $Y=750 $dt=0
M12 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=11550 $Y=750 $dt=0
M13 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=12520 $Y=750 $dt=0
M14 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=13410 $Y=750 $dt=0
M15 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=14380 $Y=750 $dt=0
M16 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.84e-13 AS=2.16e-13 PD=2.56e-06 PS=1.34e-06 $X=15270 $Y=750 $dt=0
M17 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=5.79287e-13 PD=1.86506e-06 PS=3.69506e-06 $X=475 $Y=2410 $dt=1
M18 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1315 $Y=2410 $dt=1
M19 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1865 $Y=2410 $dt=1
M20 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=2705 $Y=2410 $dt=1
M21 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=3255 $Y=2410 $dt=1
M22 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=4095 $Y=2410 $dt=1
M23 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=4645 $Y=2410 $dt=1
M24 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=5485 $Y=2410 $dt=1
M25 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=6035 $Y=2410 $dt=1
M26 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=6875 $Y=2410 $dt=1
M27 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=7425 $Y=2410 $dt=1
M28 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=8265 $Y=2410 $dt=1
M29 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=8815 $Y=2410 $dt=1
M30 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=9655 $Y=2410 $dt=1
M31 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=10205 $Y=2410 $dt=1
M32 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=11045 $Y=2410 $dt=1
M33 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=11595 $Y=2410 $dt=1
M34 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=12435 $Y=2410 $dt=1
M35 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=12985 $Y=2410 $dt=1
M36 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=13825 $Y=2410 $dt=1
M37 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=14375 $Y=2410 $dt=1
M38 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=1.15229e-12 AS=2.54913e-13 PD=4.89506e-06 PS=1.86506e-06 $X=15215 $Y=2410 $dt=1
.ends BUJI3VX16

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX0                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX0 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=4
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.923e-13 AS=2.016e-13 PD=2.005e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=3.923e-13 PD=1.8e-06 PS=2.005e-06 $X=1735 $Y=1130 $dt=0
M2 vdd3i! A 6 vdd3i! pe3i L=3e-07 W=9e-07 AD=5.7805e-13 AS=4.32e-13 PD=2.33911e-06 PS=2.76e-06 $X=620 $Y=2410 $dt=1
M3 Q 6 vdd3i! vdd3i! pe3i L=3e-07 W=1.12e-06 AD=5.376e-13 AS=7.1935e-13 PD=3.2e-06 PS=2.91089e-06 $X=1785 $Y=2410 $dt=1
.ends BUJI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA2I1JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA2I1JI3VX1 vdd3i! gnd3i! AN Q B
*.DEVICECLIMB
** N=8 EP=5 FDC=6
M0 gnd3i! AN 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.44754e-13 AS=2.016e-13 PD=1.25038e-06 PS=1.8e-06 $X=620 $Y=660 $dt=0
M1 7 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=5.18646e-13 PD=1.14e-06 PS=2.64962e-06 $X=1680 $Y=660 $dt=0
M2 Q B 7 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=1.1125e-13 PD=2.74e-06 PS=1.14e-06 $X=2280 $Y=660 $dt=0
M3 vdd3i! AN 8 vdd3i! pe3i L=3e-07 W=7e-07 AD=6.84341e-13 AS=3.36e-13 PD=3.08e-06 PS=2.36e-06 $X=620 $Y=2410 $dt=1
M4 Q 8 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.7e-13 AS=9.7763e-13 PD=1.54e-06 PS=4.4e-06 $X=1510 $Y=2410 $dt=1
M5 vdd3i! B Q vdd3i! pe3i L=3e-07 W=1e-06 AD=9.7763e-13 AS=2.7e-13 PD=4.4e-06 PS=1.54e-06 $X=2350 $Y=2410 $dt=1
.ends NA2I1JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DLY1JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DLY1JI3VX1 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=8 EP=4 FDC=8
M0 gnd3i! A 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.591e-13 AS=2.016e-13 PD=2.13e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 6 8 gnd3i! gnd3i! ne3i L=8e-07 W=4.2e-07 AD=2.415e-13 AS=3.591e-13 PD=1.99e-06 PS=2.13e-06 $X=1590 $Y=1400 $dt=0
M2 gnd3i! 6 7 gnd3i! ne3i L=1e-06 W=4.2e-07 AD=2.6662e-13 AS=2.016e-13 PD=1.28565e-06 PS=1.8e-06 $X=2860 $Y=660 $dt=0
M3 Q 7 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.3165e-13 AS=5.6498e-13 PD=2.75e-06 PS=2.72435e-06 $X=4625 $Y=660 $dt=0
M4 vdd3i! A 8 vdd3i! pe3i L=3e-07 W=6.7e-07 AD=4.61962e-13 AS=3.3835e-13 PD=2.62468e-06 PS=2.35e-06 $X=645 $Y=2680 $dt=1
M5 6 8 vdd3i! vdd3i! pe3i L=1e-06 W=4.2e-07 AD=2.00088e-13 AS=2.89588e-13 PD=1.76778e-06 PS=1.64532e-06 $X=1590 $Y=2680 $dt=1
M6 vdd3i! 6 7 vdd3i! pe3i L=7.5e-07 W=4.2e-07 AD=2.78313e-13 AS=2.00088e-13 PD=1.17049e-06 PS=1.76778e-06 $X=3110 $Y=3400 $dt=1
M7 Q 7 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.191e-13 AS=9.34337e-13 PD=3.84e-06 PS=3.92951e-06 $X=4650 $Y=2410 $dt=1
.ends DLY1JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OR4JI3VX1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OR4JI3VX1 vdd3i! gnd3i! C D Q B A
*.DEVICECLIMB
** N=13 EP=7 FDC=12
M0 11 C gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=4.12474e-13 PD=9.6e-07 PS=2.12185e-06 $X=510 $Y=1130 $dt=0
M1 gnd3i! D 11 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=4.12474e-13 AS=1.134e-13 PD=2.12185e-06 PS=9.6e-07 $X=1400 $Y=1130 $dt=0
M2 10 11 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=8.74052e-13 PD=1.14e-06 PS=4.4963e-06 $X=2330 $Y=660 $dt=0
M3 Q 9 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.56e-13 AS=1.1125e-13 PD=2.64627e-06 PS=1.14e-06 $X=2930 $Y=660 $dt=0
M4 9 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=7.908e-13 PD=9.6e-07 PS=4.27314e-06 $X=4410 $Y=1130 $dt=0
M5 gnd3i! A 9 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=7.908e-13 AS=1.134e-13 PD=4.27314e-06 PS=9.6e-07 $X=5300 $Y=1130 $dt=0
M6 13 C 11 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=4.08e-13 PD=1.1e-06 PS=2.66e-06 $X=620 $Y=2410 $dt=1
M7 vdd3i! D 13 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=6.21177e-13 AS=1.0625e-13 PD=2.08363e-06 PS=1.1e-06 $X=1170 $Y=2410 $dt=1
M8 Q 11 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=1.03042e-12 PD=1.95e-06 PS=3.45637e-06 $X=2480 $Y=2410 $dt=1
M9 vdd3i! 9 Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.09631e-12 AS=3.807e-13 PD=3.53124e-06 PS=1.95e-06 $X=3320 $Y=2410 $dt=1
M10 12 B vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=6.60894e-13 PD=1.1e-06 PS=2.12876e-06 $X=4690 $Y=2410 $dt=1
M11 9 A 12 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.08e-13 AS=1.0625e-13 PD=2.66e-06 PS=1.1e-06 $X=5240 $Y=2410 $dt=1
.ends OR4JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DFRRQJI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DFRRQJI3VX1 vdd3i! gnd3i! RN D C Q
*.DEVICECLIMB
** N=23 EP=6 FDC=30
M0 gnd3i! 17 19 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.39017e-13 AS=2.016e-13 PD=9.16947e-07 PS=1.8e-06 $X=620 $Y=660 $dt=0
M1 10 RN gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.28952e-13 AS=2.94583e-13 PD=2.36956e-06 PS=1.94305e-06 $X=1510 $Y=660 $dt=0
M2 18 19 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.55236e-13 PD=6.7e-07 PS=1.11822e-06 $X=2340 $Y=1390 $dt=0
M3 17 9 18 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=2940 $Y=1390 $dt=0
M4 16 15 17 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=3830 $Y=1390 $dt=0
M5 10 D 16 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.835e-13 AS=5.25e-14 PD=2.19e-06 PS=6.7e-07 $X=4430 $Y=1390 $dt=0
M6 gnd3i! C 15 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.659e-13 AS=2.016e-13 PD=1.21e-06 PS=1.8e-06 $X=6060 $Y=1390 $dt=0
M7 9 15 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.95e-13 AS=1.659e-13 PD=2.23e-06 PS=1.21e-06 $X=7045 $Y=1390 $dt=0
M8 14 19 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=8695 $Y=1020 $dt=0
M9 13 9 14 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=9295 $Y=1020 $dt=0
M10 12 15 13 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=10185 $Y=1020 $dt=0
M11 8 11 12 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.55817e-13 AS=5.25e-14 PD=9.68244e-07 PS=6.7e-07 $X=10785 $Y=1020 $dt=0
M12 gnd3i! RN 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=6.52289e-13 AS=3.30183e-13 PD=3.3375e-06 PS=2.05176e-06 $X=11755 $Y=660 $dt=0
M13 11 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=3.07822e-13 PD=1.8e-06 PS=1.575e-06 $X=12560 $Y=1130 $dt=0
M14 Q 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=6.52289e-13 PD=2.74e-06 PS=3.3375e-06 $X=14150 $Y=660 $dt=0
M15 vdd3i! 17 19 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=1.944e-13 AS=3.456e-13 PD=1.26e-06 PS=2.4e-06 $X=620 $Y=2670 $dt=1
M16 17 RN vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.136e-13 AS=1.944e-13 PD=2.4e-06 PS=1.26e-06 $X=1460 $Y=2670 $dt=1
M17 23 19 vdd3i! vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=5.1875e-13 PD=6.7e-07 PS=2.99e-06 $X=3080 $Y=3400 $dt=1
M18 17 15 23 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=1.21617e-13 AS=5.25e-14 PD=9.13043e-07 PS=6.7e-07 $X=3630 $Y=3400 $dt=1
M19 22 9 17 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=1.2e-13 AS=2.77983e-13 PD=1.21e-06 PS=2.08696e-06 $X=4470 $Y=2860 $dt=1
M20 vdd3i! D 22 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=5.00229e-13 AS=1.2e-13 PD=2.34286e-06 PS=1.21e-06 $X=5020 $Y=2860 $dt=1
M21 15 C vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=4.94875e-13 AS=3.75171e-13 PD=3.04e-06 PS=1.75714e-06 $X=6060 $Y=2860 $dt=1
M22 vdd3i! 15 9 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.92547e-13 AS=3.528e-13 PD=1.8586e-06 PS=2.42e-06 $X=7720 $Y=2670 $dt=1
M23 21 19 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=1.25e-13 AS=5.45203e-13 PD=1.25e-06 PS=2.5814e-06 $X=8740 $Y=2820 $dt=1
M24 13 15 21 vdd3i! pe3i L=3e-07 W=1e-06 AD=2.96338e-13 AS=1.25e-13 PD=2.19718e-06 PS=1.25e-06 $X=9290 $Y=2820 $dt=1
M25 20 9 13 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=1.24462e-13 PD=6.7e-07 PS=9.22817e-07 $X=10150 $Y=3235 $dt=1
M26 vdd3i! 11 20 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=4.10996e-13 AS=5.25e-14 PD=1.64789e-06 PS=6.7e-07 $X=10700 $Y=3235 $dt=1
M27 vdd3i! RN 13 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=7.04565e-13 AS=2.976e-13 PD=2.82495e-06 PS=2.4e-06 $X=11900 $Y=2410 $dt=1
M28 11 13 vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.456e-13 AS=7.04565e-13 PD=2.4e-06 PS=2.82495e-06 $X=12740 $Y=2410 $dt=1
M29 Q 13 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=1.37977e-12 PD=3.78e-06 PS=5.5322e-06 $X=14200 $Y=2410 $dt=1
.ends DFRRQJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INJI3VX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INJI3VX1 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=5 EP=4 FDC=2
M0 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=6e-07 AD=2.88e-13 AS=6.428e-13 PD=2.16e-06 PS=3.62e-06 $X=710 $Y=950 $dt=0
M1 Q A vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=1.0562e-12 PD=3.78e-06 PS=4.76e-06 $X=760 $Y=2410 $dt=1
.ends INJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INJI3VX2                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INJI3VX2 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=5 EP=4 FDC=4
M0 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=1.296e-13 AS=4.408e-13 PD=1.02e-06 PS=3.52e-06 $X=500 $Y=1070 $dt=0
M1 gnd3i! A Q gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=4.408e-13 AS=1.296e-13 PD=3.52e-06 PS=1.02e-06 $X=1390 $Y=1070 $dt=0
M2 Q A vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=8.151e-13 PD=1.87971e-06 PS=4.50971e-06 $X=560 $Y=2410 $dt=1
M3 vdd3i! A Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=8.01e-13 AS=2.751e-13 PD=4.48971e-06 PS=1.87971e-06 $X=1400 $Y=2410 $dt=1
.ends INJI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX12                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX12 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=28
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=4.148e-13 AS=3.84e-13 PD=1.98e-06 PS=2.56e-06 $X=620 $Y=750 $dt=0
M1 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=4.148e-13 PD=1.34e-06 PS=1.98e-06 $X=1710 $Y=750 $dt=0
M2 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=2600 $Y=750 $dt=0
M3 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=3570 $Y=750 $dt=0
M4 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=4460 $Y=750 $dt=0
M5 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=5430 $Y=750 $dt=0
M6 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=6320 $Y=750 $dt=0
M7 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=7290 $Y=750 $dt=0
M8 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=8180 $Y=750 $dt=0
M9 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=9150 $Y=750 $dt=0
M10 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.194e-13 AS=2.16e-13 PD=1.36e-06 PS=1.34e-06 $X=10040 $Y=750 $dt=0
M11 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.84e-13 AS=2.194e-13 PD=2.56e-06 PS=1.36e-06 $X=10930 $Y=750 $dt=0
M12 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=5.79287e-13 PD=1.86506e-06 PS=3.69506e-06 $X=475 $Y=2410 $dt=1
M13 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1315 $Y=2410 $dt=1
M14 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1865 $Y=2410 $dt=1
M15 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=2705 $Y=2410 $dt=1
M16 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=3255 $Y=2410 $dt=1
M17 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=4095 $Y=2410 $dt=1
M18 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=4645 $Y=2410 $dt=1
M19 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=5485 $Y=2410 $dt=1
M20 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=6035 $Y=2410 $dt=1
M21 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=6875 $Y=2410 $dt=1
M22 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=7425 $Y=2410 $dt=1
M23 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=8265 $Y=2410 $dt=1
M24 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=8815 $Y=2410 $dt=1
M25 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=9655 $Y=2410 $dt=1
M26 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=10205 $Y=2410 $dt=1
M27 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=8.53088e-13 AS=2.54913e-13 PD=4.55506e-06 PS=1.86506e-06 $X=11045 $Y=2410 $dt=1
.ends BUJI3VX12

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ON22JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ON22JI3VX1 vdd3i! gnd3i! D C Q A B
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 gnd3i! D 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=4.272e-13 PD=1.86e-06 PS=2.74e-06 $X=720 $Y=660 $dt=0
M1 9 C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=1690 $Y=660 $dt=0
M2 Q A 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=2580 $Y=660 $dt=0
M3 9 B Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.666e-13 AS=2.403e-13 PD=2.84e-06 PS=1.43e-06 $X=3470 $Y=660 $dt=0
M4 11 D vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=8.802e-13 PD=1.66e-06 PS=4.56e-06 $X=1120 $Y=2410 $dt=1
M5 Q C 11 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=1.7625e-13 PD=1.95e-06 PS=1.66e-06 $X=1670 $Y=2410 $dt=1
M6 10 A Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=3.807e-13 PD=1.66e-06 PS=1.95e-06 $X=2510 $Y=2410 $dt=1
M7 vdd3i! B 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=8.802e-13 AS=1.7625e-13 PD=4.56e-06 PS=1.66e-06 $X=3060 $Y=2410 $dt=1
.ends ON22JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AN31JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AN31JI3VX1 vdd3i! gnd3i! A B C Q D
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 10 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.335e-13 AS=6.098e-13 PD=1.19e-06 PS=3.52e-06 $X=660 $Y=660 $dt=0
M1 9 B 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.35725e-13 AS=1.335e-13 PD=1.195e-06 PS=1.19e-06 $X=1310 $Y=660 $dt=0
M2 Q C 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.0257e-13 AS=1.35725e-13 PD=1.8043e-06 PS=1.195e-06 $X=1965 $Y=660 $dt=0
M3 gnd3i! D Q gnd3i! ne3i L=3.5e-07 W=5.75e-07 AD=5.783e-13 AS=1.9548e-13 PD=3.52e-06 PS=1.1657e-06 $X=2910 $Y=975 $dt=0
M4 11 A vdd3i! vdd3i! pe3i L=3.00061e-07 W=1.44471e-06 AD=3.0525e-13 AS=5.93475e-13 PD=1.86471e-06 PS=3.72971e-06 $X=525 $Y=2425 $dt=1
M5 vdd3i! B 11 vdd3i! pe3i L=3.00061e-07 W=1.44471e-06 AD=4.42387e-13 AS=3.0525e-13 PD=2.08971e-06 PS=1.86471e-06 $X=1365 $Y=2425 $dt=1
M6 11 C vdd3i! vdd3i! pe3i L=3.00061e-07 W=1.44471e-06 AD=2.6565e-13 AS=4.42387e-13 PD=1.86471e-06 PS=2.08971e-06 $X=2310 $Y=2425 $dt=1
M7 Q D 11 vdd3i! pe3i L=3.00061e-07 W=1.44471e-06 AD=7.2375e-13 AS=2.6565e-13 PD=3.85971e-06 PS=1.86471e-06 $X=2910 $Y=2425 $dt=1
.ends AN31JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO3JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO3JI3VX0 vdd3i! gnd3i! C Q B A
*.DEVICECLIMB
** N=9 EP=6 FDC=6
M0 Q C gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.75467e-13 PD=9.6e-07 PS=2.95333e-06 $X=615 $Y=1130 $dt=0
M1 gnd3i! B Q gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.75467e-13 AS=1.134e-13 PD=2.95333e-06 PS=9.6e-07 $X=1505 $Y=1130 $dt=0
M2 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=5.75467e-13 PD=1.8e-06 PS=2.95333e-06 $X=2390 $Y=1130 $dt=0
M3 9 C vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=1.55e-13 AS=1.3584e-12 PD=1.31e-06 PS=5.15e-06 $X=955 $Y=2410 $dt=1
M4 8 B 9 vdd3i! pe3i L=3e-07 W=1e-06 AD=1.55e-13 AS=1.55e-13 PD=1.31e-06 PS=1.31e-06 $X=1565 $Y=2410 $dt=1
M5 Q A 8 vdd3i! pe3i L=3e-07 W=1e-06 AD=4.8e-13 AS=1.55e-13 PD=2.96e-06 PS=1.31e-06 $X=2175 $Y=2410 $dt=1
.ends NO3JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OR4JI3VX2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OR4JI3VX2 vdd3i! gnd3i! C D Q B A
*.DEVICECLIMB
** N=14 EP=7 FDC=16
M0 10 C gnd3i! gnd3i! ne3i L=3.5e-07 W=7e-07 AD=1.9155e-13 AS=3.417e-13 PD=1.255e-06 PS=2.39e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! D 10 gnd3i! ne3i L=3.5e-07 W=7e-07 AD=2.07711e-13 AS=1.9155e-13 PD=1.27673e-06 PS=1.255e-06 $X=1510 $Y=660 $dt=0
M2 12 10 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=2.64089e-13 PD=1.14e-06 PS=1.62327e-06 $X=2420 $Y=660 $dt=0
M3 Q 9 12 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=1.1125e-13 PD=1.43e-06 PS=1.14e-06 $X=3020 $Y=660 $dt=0
M4 11 9 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.2015e-13 AS=2.403e-13 PD=1.16e-06 PS=1.43e-06 $X=3910 $Y=660 $dt=0
M5 gnd3i! 10 11 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.54126e-13 AS=1.2015e-13 PD=1.60088e-06 PS=1.16e-06 $X=4530 $Y=660 $dt=0
M6 9 B gnd3i! gnd3i! ne3i L=3.5e-07 W=7e-07 AD=1.9155e-13 AS=1.99874e-13 PD=1.255e-06 PS=1.25912e-06 $X=5420 $Y=660 $dt=0
M7 gnd3i! A 9 gnd3i! ne3i L=3.5e-07 W=7e-07 AD=3.417e-13 AS=1.9155e-13 PD=2.39e-06 PS=1.255e-06 $X=6310 $Y=660 $dt=0
M8 14 C 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=6.768e-13 PD=1.66e-06 PS=3.78e-06 $X=710 $Y=2410 $dt=1
M9 vdd3i! D 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=5.47043e-13 AS=1.7625e-13 PD=2.41704e-06 PS=1.66e-06 $X=1260 $Y=2410 $dt=1
M10 Q 10 vdd3i! vdd3i! pe3i L=2.99799e-07 W=1.41828e-06 AD=3.622e-13 AS=5.50257e-13 PD=1.93828e-06 PS=2.43124e-06 $X=2210 $Y=2410 $dt=1
M11 vdd3i! 9 Q vdd3i! pe3i L=2.99799e-07 W=1.41828e-06 AD=4.987e-13 AS=3.622e-13 PD=2.36828e-06 PS=1.93828e-06 $X=3050 $Y=2410 $dt=1
M12 Q 9 vdd3i! vdd3i! pe3i L=2.99799e-07 W=1.41828e-06 AD=3.622e-13 AS=4.987e-13 PD=1.93828e-06 PS=2.36828e-06 $X=3930 $Y=2410 $dt=1
M13 vdd3i! 10 Q vdd3i! pe3i L=2.99799e-07 W=1.41828e-06 AD=5.8556e-13 AS=3.622e-13 PD=2.47136e-06 PS=1.93828e-06 $X=4770 $Y=2410 $dt=1
M14 13 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=5.8214e-13 PD=1.66e-06 PS=2.45692e-06 $X=5760 $Y=2410 $dt=1
M15 9 A 13 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=1.7625e-13 PD=3.78e-06 PS=1.66e-06 $X=6310 $Y=2410 $dt=1
.ends OR4JI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: HAJI3VX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt HAJI3VX1 vdd3i! gnd3i! S B A CO
*.DEVICECLIMB
** N=12 EP=6 FDC=14
M0 gnd3i! 8 S gnd3i! ne3i L=3.49889e-07 W=8.98284e-07 AD=4.998e-13 AS=4.174e-13 PD=3.41456e-06 PS=2.72828e-06 $X=600 $Y=660 $dt=0
M1 gnd3i! A 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.52e-13 PD=1.43e-06 PS=2.74e-06 $X=2070 $Y=660 $dt=0
M2 9 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.70969e-13 AS=2.403e-13 PD=1.71986e-06 PS=1.43e-06 $X=2960 $Y=660 $dt=0
M3 8 10 9 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=3.632e-13 AS=1.79631e-13 PD=2.84284e-06 PS=1.14014e-06 $X=3850 $Y=960 $dt=0
M4 gnd3i! 10 CO gnd3i! ne3i L=3.5e-07 W=5.5e-07 AD=1.56292e-13 AS=2.4195e-13 PD=1.09236e-06 PS=2.03071e-06 $X=5380 $Y=1000 $dt=0
M5 11 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=2.52908e-13 PD=1.14e-06 PS=1.76764e-06 $X=6270 $Y=660 $dt=0
M6 10 A 11 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=1.1125e-13 PD=2.74e-06 PS=1.14e-06 $X=6870 $Y=660 $dt=0
M7 vdd3i! 8 S vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.07833e-13 AS=7.1205e-13 PD=2.97939e-06 PS=3.83e-06 $X=645 $Y=2410 $dt=1
M8 12 A vdd3i! vdd3i! pe3i L=3e-07 W=8.9e-07 AD=1.335e-13 AS=3.83667e-13 PD=1.19e-06 PS=1.88061e-06 $X=1615 $Y=2630 $dt=1
M9 8 B 12 vdd3i! pe3i L=3e-07 W=8.9e-07 AD=4.9565e-13 AS=1.335e-13 PD=2.12e-06 PS=1.19e-06 $X=2215 $Y=2630 $dt=1
M10 vdd3i! 10 8 vdd3i! pe3i L=3e-07 W=8.9e-07 AD=4.8925e-13 AS=4.9565e-13 PD=3.49e-06 PS=2.12e-06 $X=3525 $Y=2630 $dt=1
M11 vdd3i! 10 CO vdd3i! pe3i L=3e-07 W=1.11e-06 AD=4.3695e-13 AS=4.7415e-13 PD=2.09e-06 PS=3.23e-06 $X=4995 $Y=2410 $dt=1
M12 10 B vdd3i! vdd3i! pe3i L=3e-07 W=1.11e-06 AD=3.2745e-13 AS=4.3695e-13 PD=1.7e-06 PS=2.09e-06 $X=5965 $Y=2410 $dt=1
M13 vdd3i! A 10 vdd3i! pe3i L=3e-07 W=1.11e-06 AD=8.7795e-13 AS=3.2745e-13 PD=4.61e-06 PS=1.7e-06 $X=6855 $Y=2410 $dt=1
.ends HAJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DLY4JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DLY4JI3VX1 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=12 EP=4 FDC=12
M0 gnd3i! A 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.323e-13 AS=2.016e-13 PD=1.05e-06 PS=1.8e-06 $X=620 $Y=660 $dt=0
M1 8 10 gnd3i! gnd3i! ne3i L=1.8e-06 W=4.2e-07 AD=1.736e-13 AS=1.323e-13 PD=1.58e-06 PS=1.05e-06 $X=1600 $Y=660 $dt=0
M2 8 10 9 gnd3i! ne3i L=1.8e-06 W=4.2e-07 AD=1.736e-13 AS=2.00088e-13 PD=1.58e-06 PS=1.76778e-06 $X=1600 $Y=1360 $dt=0
M3 gnd3i! 9 7 gnd3i! ne3i L=1.1e-06 W=4.2e-07 AD=4.30324e-13 AS=2.16e-13 PD=1.75053e-06 PS=1.66e-06 $X=4630 $Y=660 $dt=0
M4 6 9 7 gnd3i! ne3i L=1.1e-06 W=4.2e-07 AD=2.00088e-13 AS=2.16e-13 PD=1.76778e-06 PS=1.66e-06 $X=4630 $Y=1400 $dt=0
M5 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.4055e-13 AS=9.11876e-13 PD=2.77e-06 PS=3.70947e-06 $X=7220 $Y=660 $dt=0
M6 vdd3i! A 10 vdd3i! pe3i L=3e-07 W=7e-07 AD=5.26875e-13 AS=3.535e-13 PD=3.30625e-06 PS=2.41e-06 $X=645 $Y=2680 $dt=1
M7 12 10 9 vdd3i! pe3i L=1.2e-06 W=4.2e-07 AD=1.674e-13 AS=2.016e-13 PD=1.56e-06 PS=1.8e-06 $X=2100 $Y=2680 $dt=1
M8 12 10 vdd3i! vdd3i! pe3i L=1.2e-06 W=4.2e-07 AD=1.674e-13 AS=3.16125e-13 PD=1.56e-06 PS=1.98375e-06 $X=2100 $Y=3400 $dt=1
M9 6 9 11 vdd3i! pe3i L=1.9e-06 W=4.2e-07 AD=2.016e-13 AS=1.674e-13 PD=1.8e-06 PS=1.56e-06 $X=4220 $Y=2680 $dt=1
M10 vdd3i! 9 11 vdd3i! pe3i L=1.9e-06 W=4.2e-07 AD=2.6367e-13 AS=1.674e-13 PD=1.32426e-06 PS=1.56e-06 $X=4220 $Y=3400 $dt=1
M11 Q 6 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.332e-13 AS=8.8518e-13 PD=3.86e-06 PS=4.44574e-06 $X=7245 $Y=2410 $dt=1
.ends DLY4JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO2I1JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO2I1JI3VX1 vdd3i! gnd3i! AN Q B
*.DEVICECLIMB
** N=8 EP=5 FDC=6
M0 gnd3i! AN 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.78131e-13 AS=2.016e-13 PD=1.19267e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 Q 7 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.4285e-13 AS=3.77469e-13 PD=1.445e-06 PS=2.52733e-06 $X=1460 $Y=660 $dt=0
M2 gnd3i! B Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=6.098e-13 AS=2.4285e-13 PD=3.52e-06 PS=1.445e-06 $X=2350 $Y=660 $dt=0
M3 vdd3i! AN 7 vdd3i! pe3i L=3e-07 W=7e-07 AD=4.32009e-13 AS=3.36e-13 PD=1.71185e-06 PS=2.36e-06 $X=620 $Y=2410 $dt=1
M4 8 7 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=8.70191e-13 PD=1.66e-06 PS=3.44815e-06 $X=1740 $Y=2410 $dt=1
M5 Q B 8 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=1.7625e-13 PD=3.78e-06 PS=1.66e-06 $X=2290 $Y=2410 $dt=1
.ends NO2I1JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AO22JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AO22JI3VX1 vdd3i! gnd3i! B A C D Q
*.DEVICECLIMB
** N=12 EP=7 FDC=10
M0 11 B gnd3i! gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=5.768e-13 PD=8.1e-07 PS=3.52e-06 $X=660 $Y=990 $dt=0
M1 10 A 11 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=1.68e-13 AS=7e-14 PD=1.16e-06 PS=8.1e-07 $X=1260 $Y=990 $dt=0
M2 9 C 10 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=1.68e-13 PD=8.1e-07 PS=1.16e-06 $X=2210 $Y=990 $dt=0
M3 gnd3i! D 9 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=3.96017e-13 AS=7e-14 PD=1.66069e-06 PS=8.1e-07 $X=2810 $Y=990 $dt=0
M4 Q 10 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=6.29383e-13 PD=2.74e-06 PS=2.63931e-06 $X=4070 $Y=660 $dt=0
M5 vdd3i! B 12 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=2.295e-13 AS=4.868e-13 PD=1.39e-06 PS=3.75e-06 $X=460 $Y=2490 $dt=1
M6 12 A vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.868e-13 AS=2.295e-13 PD=3.75e-06 PS=1.39e-06 $X=1300 $Y=2490 $dt=1
M7 10 C 12 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=2.295e-13 AS=4.868e-13 PD=1.39e-06 PS=3.75e-06 $X=2020 $Y=2490 $dt=1
M8 12 D 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.868e-13 AS=2.295e-13 PD=3.75e-06 PS=1.39e-06 $X=2860 $Y=2490 $dt=1
M9 Q 10 vdd3i! vdd3i! pe3i L=3.01705e-07 W=1.47627e-06 AD=5.312e-13 AS=7.778e-13 PD=3.68627e-06 PS=4.46627e-06 $X=4120 $Y=2410 $dt=1
.ends AO22JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX6                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX6 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=14
M0 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=6.008e-13 PD=1.34e-06 PS=3.52e-06 $X=660 $Y=750 $dt=0
M1 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=5.84805e-13 AS=2.16e-13 PD=2.17751e-06 PS=1.34e-06 $X=1550 $Y=750 $dt=0
M2 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=6.50595e-13 PD=1.43e-06 PS=2.42249e-06 $X=2960 $Y=660 $dt=0
M3 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=3850 $Y=660 $dt=0
M4 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=4820 $Y=660 $dt=0
M5 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=6.098e-13 AS=2.403e-13 PD=3.52e-06 PS=1.43e-06 $X=5710 $Y=660 $dt=0
M6 6 A vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=6.3285e-13 PD=1.87971e-06 PS=3.75971e-06 $X=525 $Y=2410 $dt=1
M7 vdd3i! A 6 vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=3.7905e-13 AS=2.751e-13 PD=1.98971e-06 PS=1.87971e-06 $X=1365 $Y=2410 $dt=1
M8 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=3.7905e-13 PD=1.87971e-06 PS=1.98971e-06 $X=2075 $Y=2410 $dt=1
M9 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=3.3675e-13 AS=2.751e-13 PD=1.92971e-06 PS=1.87971e-06 $X=2915 $Y=2410 $dt=1
M10 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=3.3675e-13 PD=1.87971e-06 PS=1.92971e-06 $X=3565 $Y=2410 $dt=1
M11 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=3.3675e-13 AS=2.751e-13 PD=1.92971e-06 PS=1.87971e-06 $X=4405 $Y=2410 $dt=1
M12 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=3.3675e-13 PD=1.87971e-06 PS=1.92971e-06 $X=5055 $Y=2410 $dt=1
M13 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=6.3285e-13 AS=2.751e-13 PD=3.75971e-06 PS=1.87971e-06 $X=5895 $Y=2410 $dt=1
.ends BUJI3VX6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ON31JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ON31JI3VX1 vdd3i! gnd3i! A B C Q D
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 9 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=6.098e-13 PD=1.43e-06 PS=3.52e-06 $X=660 $Y=660 $dt=0
M1 gnd3i! B 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=1550 $Y=660 $dt=0
M2 9 C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=2520 $Y=660 $dt=0
M3 Q D 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=2.403e-13 PD=2.74e-06 PS=1.43e-06 $X=3410 $Y=660 $dt=0
M4 11 A vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=9.066e-13 PD=1.72e-06 PS=4.59e-06 $X=1145 $Y=2410 $dt=1
M5 10 B 11 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=2.1855e-13 PD=1.72e-06 PS=1.72e-06 $X=1755 $Y=2410 $dt=1
M6 Q C 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=5.30442e-13 AS=2.1855e-13 PD=2.60067e-06 PS=1.72e-06 $X=2365 $Y=2410 $dt=1
M7 vdd3i! D Q vdd3i! pe3i L=3e-07 W=8.4e-07 AD=1.1576e-12 AS=3.16008e-13 PD=4.94e-06 PS=1.54933e-06 $X=3330 $Y=2410 $dt=1
.ends ON31JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: EO3JI3VX1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt EO3JI3VX1 vdd3i! gnd3i! C B A Q
*.DEVICECLIMB
** N=16 EP=6 FDC=20
M0 12 C gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.628e-13 PD=9.6e-07 PS=3.52e-06 $X=660 $Y=1130 $dt=0
M1 gnd3i! B 12 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.30196e-13 AS=1.134e-13 PD=1.36723e-06 PS=9.6e-07 $X=1550 $Y=1130 $dt=0
M2 11 C gnd3i! gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=6.5e-14 AS=2.85004e-13 PD=7.7e-07 PS=1.69277e-06 $X=2910 $Y=1030 $dt=0
M3 10 B 11 gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=1.404e-13 AS=6.5e-14 PD=1.06e-06 PS=7.7e-07 $X=3510 $Y=1030 $dt=0
M4 gnd3i! 12 10 gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=8.05779e-13 AS=1.404e-13 PD=2.83787e-06 PS=1.06e-06 $X=4400 $Y=1030 $dt=0
M5 9 10 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=6.50821e-13 PD=9.6e-07 PS=2.29213e-06 $X=6075 $Y=1130 $dt=0
M6 gnd3i! A 9 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.90537e-13 AS=1.134e-13 PD=1.53255e-06 PS=9.6e-07 $X=6965 $Y=1130 $dt=0
M7 8 A gnd3i! gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=6.5e-14 AS=3.59713e-13 PD=7.7e-07 PS=1.89745e-06 $X=8140 $Y=1030 $dt=0
M8 Q 10 8 gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=1.404e-13 AS=6.5e-14 PD=1.06e-06 PS=7.7e-07 $X=8740 $Y=1030 $dt=0
M9 gnd3i! 9 Q gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=5.728e-13 AS=1.404e-13 PD=3.52e-06 PS=1.06e-06 $X=9630 $Y=1030 $dt=0
M10 16 C vdd3i! vdd3i! pe3i L=3e-07 W=1.3e-06 AD=1.95e-13 AS=6.603e-13 PD=1.6e-06 PS=3.63e-06 $X=645 $Y=2520 $dt=1
M11 12 B 16 vdd3i! pe3i L=3e-07 W=1.3e-06 AD=5.157e-13 AS=1.95e-13 PD=3.61e-06 PS=1.6e-06 $X=1245 $Y=2520 $dt=1
M12 vdd3i! C 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=5.8645e-13 PD=2e-06 PS=3.83e-06 $X=2675 $Y=2410 $dt=1
M13 14 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=4.1595e-13 PD=2e-06 PS=2e-06 $X=3565 $Y=2410 $dt=1
M14 10 12 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=5.6965e-13 AS=4.1595e-13 PD=3.83e-06 PS=2e-06 $X=4455 $Y=2410 $dt=1
M15 15 10 vdd3i! vdd3i! pe3i L=3e-07 W=1.3e-06 AD=1.95e-13 AS=5.301e-13 PD=1.6e-06 PS=3.61e-06 $X=5885 $Y=2410 $dt=1
M16 9 A 15 vdd3i! pe3i L=3e-07 W=1.3e-06 AD=5.157e-13 AS=1.95e-13 PD=3.61e-06 PS=1.6e-06 $X=6485 $Y=2410 $dt=1
M17 vdd3i! A 13 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=5.8645e-13 PD=2e-06 PS=3.83e-06 $X=7915 $Y=2410 $dt=1
M18 13 10 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=4.1595e-13 PD=2e-06 PS=2e-06 $X=8805 $Y=2410 $dt=1
M19 Q 9 13 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.1205e-13 AS=4.1595e-13 PD=3.83e-06 PS=2e-06 $X=9695 $Y=2410 $dt=1
.ends EO3JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX2                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX2 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=6
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=6e-07 AD=2.96727e-13 AS=2.88e-13 PD=1.69091e-06 PS=2.16e-06 $X=620 $Y=950 $dt=0
M1 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=7.2e-07 AD=2.016e-13 AS=3.56073e-13 PD=1.512e-06 PS=2.02909e-06 $X=1590 $Y=830 $dt=0
M2 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=4.648e-13 AS=1.344e-13 PD=3.52e-06 PS=1.008e-06 $X=2480 $Y=1070 $dt=0
M3 vdd3i! A 6 vdd3i! pe3i L=3e-07 W=1.1e-06 AD=5.39943e-13 AS=5.28e-13 PD=2.20442e-06 PS=3.16e-06 $X=620 $Y=2410 $dt=1
M4 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=7.16507e-13 PD=1.87971e-06 PS=2.92528e-06 $X=1640 $Y=2410 $dt=1
M5 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=8.6265e-13 AS=2.751e-13 PD=4.56971e-06 PS=1.87971e-06 $X=2480 $Y=2410 $dt=1
.ends BUJI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INJI3VX3                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INJI3VX3 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=5 EP=4 FDC=5
M0 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=7.586e-13 PD=1.43e-06 PS=3.76e-06 $X=780 $Y=660 $dt=0
M1 gnd3i! A Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=7.586e-13 AS=2.403e-13 PD=3.76e-06 PS=1.43e-06 $X=1670 $Y=660 $dt=0
M2 Q A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=6.12287e-13 PD=1.86506e-06 PS=3.78506e-06 $X=490 $Y=2410 $dt=1
M3 vdd3i! A Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.86587e-13 AS=2.54913e-13 PD=1.88506e-06 PS=1.86506e-06 $X=1330 $Y=2410 $dt=1
M4 Q A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=5.51013e-13 AS=2.86587e-13 PD=3.69506e-06 PS=1.88506e-06 $X=1880 $Y=2410 $dt=1
.ends INJI3VX3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA3I2JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA3I2JI3VX1 vdd3i! gnd3i! AN BN C Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 9 AN gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=4.00432e-13 PD=9.6e-07 PS=2.10243e-06 $X=540 $Y=1130 $dt=0
M1 gnd3i! BN 9 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=4.00432e-13 AS=1.134e-13 PD=2.10243e-06 PS=9.6e-07 $X=1430 $Y=1130 $dt=0
M2 8 C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=8.48535e-13 PD=1.14e-06 PS=4.45514e-06 $X=2290 $Y=660 $dt=0
M3 Q 9 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.806e-13 AS=1.1125e-13 PD=2.86e-06 PS=1.14e-06 $X=2890 $Y=660 $dt=0
M4 10 AN 9 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=4.08e-13 PD=1.1e-06 PS=2.66e-06 $X=620 $Y=2410 $dt=1
M5 vdd3i! BN 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=7.38476e-13 AS=1.0625e-13 PD=3.31526e-06 PS=1.1e-06 $X=1170 $Y=2410 $dt=1
M6 vdd3i! C Q vdd3i! pe3i L=3.00037e-07 W=1.00071e-06 AD=8.69412e-13 AS=2.376e-13 PD=3.90308e-06 PS=1.49071e-06 $X=2170 $Y=2410 $dt=1
M7 Q 9 vdd3i! vdd3i! pe3i L=3.00037e-07 W=1.00071e-06 AD=2.376e-13 AS=8.69412e-13 PD=1.49071e-06 PS=3.90308e-06 $X=3010 $Y=2410 $dt=1
.ends NA3I2JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: EN3JI3VX1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt EN3JI3VX1 vdd3i! gnd3i! C B A Q
*.DEVICECLIMB
** N=16 EP=6 FDC=20
M0 13 C gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=2.016e-13 PD=9.6e-07 PS=1.8e-06 $X=620 $Y=1030 $dt=0
M1 gnd3i! B 13 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.97668e-13 AS=1.134e-13 PD=1.24213e-06 PS=9.6e-07 $X=1510 $Y=1030 $dt=0
M2 12 C gnd3i! gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=6.5e-14 AS=2.44732e-13 PD=7.7e-07 PS=1.53787e-06 $X=2730 $Y=930 $dt=0
M3 11 B 12 gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=1.404e-13 AS=6.5e-14 PD=1.06e-06 PS=7.7e-07 $X=3330 $Y=930 $dt=0
M4 gnd3i! 13 11 gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=5.308e-13 AS=1.404e-13 PD=3.32e-06 PS=1.06e-06 $X=4220 $Y=930 $dt=0
M5 9 11 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=5850 $Y=970 $dt=0
M6 gnd3i! A 9 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=6450 $Y=970 $dt=0
M7 8 A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=1.134e-13 PD=9.6e-07 PS=9.6e-07 $X=7340 $Y=970 $dt=0
M8 gnd3i! 11 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.965e-13 AS=1.134e-13 PD=3.17071e-06 PS=9.6e-07 $X=8230 $Y=970 $dt=0
M9 Q 10 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=2.0035e-13 PD=1.8e-06 PS=1.77071e-06 $X=9670 $Y=1130 $dt=0
M10 16 C vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.115e-13 AS=7.1585e-13 PD=1.71e-06 PS=3.85e-06 $X=645 $Y=2410 $dt=1
M11 13 B 16 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=5.5365e-13 AS=2.115e-13 PD=3.83e-06 PS=1.71e-06 $X=1245 $Y=2410 $dt=1
M12 vdd3i! C 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.23e-13 AS=5.8645e-13 PD=2.01e-06 PS=3.83e-06 $X=2675 $Y=2410 $dt=1
M13 14 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=4.23e-13 PD=2e-06 PS=2.01e-06 $X=3575 $Y=2410 $dt=1
M14 11 13 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.1205e-13 AS=4.1595e-13 PD=3.83e-06 PS=2e-06 $X=4465 $Y=2410 $dt=1
M15 10 11 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=9.1545e-13 PD=2e-06 PS=4.61e-06 $X=6095 $Y=2410 $dt=1
M16 vdd3i! A 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.956e-13 AS=4.1595e-13 PD=2.63e-06 PS=2e-06 $X=6985 $Y=2410 $dt=1
M17 15 A vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.115e-13 AS=6.956e-13 PD=1.71e-06 PS=2.63e-06 $X=8155 $Y=2410 $dt=1
M18 Q 11 15 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.66787e-13 AS=2.115e-13 PD=2.36668e-06 PS=1.71e-06 $X=8755 $Y=2410 $dt=1
M19 vdd3i! 10 Q vdd3i! pe3i L=3e-07 W=9.85e-07 AD=8.62325e-13 AS=3.26088e-13 PD=4.61e-06 PS=1.65332e-06 $X=9655 $Y=2410 $dt=1
.ends EN3JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: SDFRRQJI3VX1                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt SDFRRQJI3VX1 vdd3i! gnd3i! SE SD RN D C Q
*.DEVICECLIMB
** N=31 EP=8 FDC=39
M0 gnd3i! SE 25 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.11575e-13 AS=2.016e-13 PD=1.6275e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 13 RN gnd3i! gnd3i! ne3i L=3.5e-07 W=5.4e-07 AD=2.079e-13 AS=2.72025e-13 PD=1.4625e-06 PS=2.0925e-06 $X=1410 $Y=660 $dt=0
M2 24 SE 13 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.617e-13 PD=6.7e-07 PS=1.1375e-06 $X=2340 $Y=960 $dt=0
M3 12 SD 24 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.163e-13 AS=5.25e-14 PD=1.45e-06 PS=6.7e-07 $X=2940 $Y=960 $dt=0
M4 23 D 12 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.163e-13 PD=6.7e-07 PS=1.45e-06 $X=3910 $Y=1000 $dt=0
M5 13 25 23 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=5.25e-14 PD=1.8e-06 PS=6.7e-07 $X=4510 $Y=1000 $dt=0
M6 gnd3i! 20 22 gnd3i! ne3i L=3.5e-07 W=7.2e-07 AD=3.01862e-13 AS=3.456e-13 PD=1.65084e-06 PS=2.4e-06 $X=6100 $Y=1090 $dt=0
M7 11 RN gnd3i! gnd3i! ne3i L=3.5e-07 W=8.85e-07 AD=2.20538e-13 AS=3.71038e-13 PD=1.77e-06 PS=2.02916e-06 $X=7070 $Y=925 $dt=0
M8 21 22 11 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.04662e-13 PD=6.7e-07 PS=8.4e-07 $X=7840 $Y=1390 $dt=0
M9 20 18 21 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=8440 $Y=1390 $dt=0
M10 12 19 20 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=1.134e-13 PD=1.8e-06 PS=9.6e-07 $X=9330 $Y=1390 $dt=0
M11 gnd3i! C 19 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.722e-13 AS=2.016e-13 PD=1.24e-06 PS=1.8e-06 $X=10920 $Y=1390 $dt=0
M12 18 19 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=1.722e-13 PD=1.8e-06 PS=1.24e-06 $X=11930 $Y=1390 $dt=0
M13 17 22 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=13520 $Y=1020 $dt=0
M14 16 18 17 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=14120 $Y=1020 $dt=0
M15 15 19 16 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=15010 $Y=1020 $dt=0
M16 10 14 15 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.47785e-13 AS=5.25e-14 PD=9.42595e-07 PS=6.7e-07 $X=15610 $Y=1020 $dt=0
M17 gnd3i! RN 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.9815e-13 AS=3.13165e-13 PD=1.56e-06 PS=1.9974e-06 $X=16540 $Y=660 $dt=0
M18 14 16 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=2.9815e-13 PD=2.74e-06 PS=1.56e-06 $X=17560 $Y=660 $dt=0
M19 Q 16 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=6.098e-13 PD=2.74e-06 PS=3.52e-06 $X=19190 $Y=660 $dt=0
M20 vdd3i! SE 25 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=5.776e-13 AS=3.456e-13 PD=2.10667e-06 PS=2.4e-06 $X=620 $Y=2800 $dt=1
M21 31 25 vdd3i! vdd3i! pe3i L=3e-07 W=9e-07 AD=1.125e-13 AS=7.22e-13 PD=1.15e-06 PS=2.63333e-06 $X=2030 $Y=2620 $dt=1
M22 28 SD 31 vdd3i! pe3i L=3e-07 W=9e-07 AD=2.43e-13 AS=1.125e-13 PD=1.44e-06 PS=1.15e-06 $X=2580 $Y=2620 $dt=1
M23 30 D 28 vdd3i! pe3i L=3e-07 W=9e-07 AD=1.125e-13 AS=2.43e-13 PD=1.15e-06 PS=1.44e-06 $X=3420 $Y=2620 $dt=1
M24 vdd3i! SE 30 vdd3i! pe3i L=3e-07 W=9e-07 AD=3.80558e-13 AS=1.125e-13 PD=1.98274e-06 PS=1.15e-06 $X=3970 $Y=2620 $dt=1
M25 22 20 vdd3i! vdd3i! pe3i L=3e-07 W=1.07e-06 AD=5.136e-13 AS=4.52442e-13 PD=3.1e-06 PS=2.35726e-06 $X=4890 $Y=2745 $dt=1
M26 vdd3i! RN 20 vdd3i! pe3i L=3e-07 W=1.02e-06 AD=9.30148e-13 AS=4.896e-13 PD=3.58417e-06 PS=3e-06 $X=6430 $Y=2800 $dt=1
M27 29 22 vdd3i! vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=3.83002e-13 PD=6.7e-07 PS=1.47583e-06 $X=7890 $Y=3060 $dt=1
M28 20 19 29 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=1.218e-13 AS=5.25e-14 PD=9.22677e-07 PS=6.7e-07 $X=8440 $Y=3060 $dt=1
M29 28 18 20 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.08e-13 AS=2.465e-13 PD=2.66e-06 PS=1.86732e-06 $X=9285 $Y=2670 $dt=1
M30 19 C vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.0675e-13 AS=6.327e-13 PD=2.37071e-06 PS=3.56e-06 $X=10970 $Y=2735 $dt=1
M31 vdd3i! 19 18 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.27981e-13 AS=4.01587e-13 PD=1.59258e-06 PS=3.03778e-06 $X=12390 $Y=2800 $dt=1
M32 27 22 vdd3i! vdd3i! pe3i L=3e-07 W=7.9e-07 AD=1.16525e-13 AS=3.59869e-13 PD=1.085e-06 PS=1.74742e-06 $X=13570 $Y=2730 $dt=1
M33 16 19 27 vdd3i! pe3i L=3e-07 W=7.9e-07 AD=2.25379e-13 AS=1.16525e-13 PD=1.73669e-06 PS=1.085e-06 $X=14165 $Y=2730 $dt=1
M34 26 18 16 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=1.19821e-13 PD=6.7e-07 PS=9.23306e-07 $X=15005 $Y=3100 $dt=1
M35 vdd3i! 14 26 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=6.29844e-13 AS=5.25e-14 PD=2.86017e-06 PS=6.7e-07 $X=15555 $Y=3100 $dt=1
M36 vdd3i! RN 16 vdd3i! pe3i L=3e-07 W=7.9e-07 AD=1.18471e-12 AS=3.19387e-13 PD=5.37983e-06 PS=2.5195e-06 $X=16775 $Y=2410 $dt=1
M37 vdd3i! 16 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=6.768e-13 PD=1.95e-06 PS=3.78e-06 $X=18400 $Y=2410 $dt=1
M38 Q 16 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=3.807e-13 PD=3.78e-06 PS=1.95e-06 $X=19240 $Y=2410 $dt=1
.ends SDFRRQJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO2JI3VX0 vdd3i! gnd3i! B Q A
*.DEVICECLIMB
** N=7 EP=5 FDC=4
M0 Q B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=7.244e-13 PD=9.6e-07 PS=4.14e-06 $X=500 $Y=1130 $dt=0
M1 gnd3i! A Q gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=7.244e-13 AS=1.134e-13 PD=4.14e-06 PS=9.6e-07 $X=1390 $Y=1130 $dt=0
M2 7 B vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=9.298e-13 PD=1.1e-06 PS=4.68e-06 $X=720 $Y=2410 $dt=1
M3 Q A 7 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.08e-13 AS=1.0625e-13 PD=2.66e-06 PS=1.1e-06 $X=1270 $Y=2410 $dt=1
.ends NO2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA4JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA4JI3VX0 vdd3i! gnd3i! D Q C B A
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 11 D gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=1.2e-13 AS=7.868e-13 PD=1.1e-06 PS=3.82e-06 $X=810 $Y=750 $dt=0
M1 10 C 11 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=1.2e-13 AS=1.2e-13 PD=1.1e-06 PS=1.1e-06 $X=1460 $Y=750 $dt=0
M2 9 B 10 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=1.2e-13 AS=1.2e-13 PD=1.1e-06 PS=1.1e-06 $X=2110 $Y=750 $dt=0
M3 Q A 9 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.84e-13 AS=1.2e-13 PD=2.56e-06 PS=1.1e-06 $X=2760 $Y=750 $dt=0
M4 Q D vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=9.882e-13 PD=1.24e-06 PS=3.92e-06 $X=540 $Y=2410 $dt=1
M5 vdd3i! C Q vdd3i! pe3i L=3e-07 W=7e-07 AD=9.882e-13 AS=1.89e-13 PD=3.92e-06 PS=1.24e-06 $X=1380 $Y=2410 $dt=1
M6 Q B vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=9.882e-13 PD=1.24e-06 PS=3.92e-06 $X=2240 $Y=2410 $dt=1
M7 vdd3i! A Q vdd3i! pe3i L=3e-07 W=7e-07 AD=9.882e-13 AS=1.89e-13 PD=3.92e-06 PS=1.24e-06 $X=3080 $Y=2410 $dt=1
.ends NA4JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA2JI3VX0 vdd3i! gnd3i! B Q A
*.DEVICECLIMB
** N=7 EP=5 FDC=4
M0 7 B gnd3i! gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=5.892e-13 PD=8.1e-07 PS=3.54e-06 $X=670 $Y=990 $dt=0
M1 Q A 7 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=2.688e-13 AS=7e-14 PD=2.08e-06 PS=8.1e-07 $X=1270 $Y=990 $dt=0
M2 Q B vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=1.1114e-12 PD=1.24e-06 PS=4.94e-06 $X=550 $Y=2410 $dt=1
M3 vdd3i! A Q vdd3i! pe3i L=3e-07 W=7e-07 AD=1.1114e-12 AS=1.89e-13 PD=4.94e-06 PS=1.24e-06 $X=1390 $Y=2410 $dt=1
.ends NA2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ON21JI3VX4                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ON21JI3VX4 vdd3i! gnd3i! B A C Q
*.DEVICECLIMB
** N=11 EP=6 FDC=16
M0 gnd3i! B 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=4.272e-13 PD=1.43e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 10 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=1510 $Y=660 $dt=0
M2 9 C 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.868e-13 AS=2.403e-13 PD=2.70971e-06 PS=1.43e-06 $X=2400 $Y=660 $dt=0
M3 gnd3i! 9 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.35783e-13 AS=4.34e-13 PD=1.42065e-06 PS=2.92971e-06 $X=3930 $Y=660 $dt=0
M4 Q 8 gnd3i! gnd3i! ne3i L=3.49164e-07 W=8.96213e-07 AD=2.32912e-13 AS=2.37429e-13 PD=1.42121e-06 PS=1.43057e-06 $X=4820 $Y=660 $dt=0
M5 gnd3i! 8 Q gnd3i! ne3i L=3.49164e-07 W=8.96213e-07 AD=2.32912e-13 AS=2.32912e-13 PD=1.42121e-06 PS=1.42121e-06 $X=5680 $Y=660 $dt=0
M6 Q 8 gnd3i! gnd3i! ne3i L=3.49164e-07 W=8.96213e-07 AD=2.32912e-13 AS=2.32912e-13 PD=1.42121e-06 PS=1.42121e-06 $X=6570 $Y=660 $dt=0
M7 gnd3i! 8 Q gnd3i! ne3i L=3.49164e-07 W=8.96213e-07 AD=4.19812e-13 AS=2.32912e-13 PD=2.73121e-06 PS=1.42121e-06 $X=7430 $Y=660 $dt=0
M8 11 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=9.418e-13 PD=1.66e-06 PS=4.63e-06 $X=695 $Y=2410 $dt=1
M9 9 A 11 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.68825e-13 AS=1.7625e-13 PD=2.075e-06 PS=1.66e-06 $X=1245 $Y=2410 $dt=1
M10 vdd3i! C 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.285e-12 AS=4.68825e-13 PD=5.02e-06 PS=2.075e-06 $X=2210 $Y=2410 $dt=1
M11 vdd3i! 9 8 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=5.48179e-13 AS=6.768e-13 PD=2.4141e-06 PS=3.78e-06 $X=4020 $Y=2410 $dt=1
M12 Q 8 vdd3i! vdd3i! pe3i L=3.00021e-07 W=1.42657e-06 AD=3.433e-13 AS=5.54621e-13 PD=1.92657e-06 PS=2.44247e-06 $X=4960 $Y=2410 $dt=1
M13 vdd3i! 8 Q vdd3i! pe3i L=3.00021e-07 W=1.42657e-06 AD=4.866e-13 AS=3.433e-13 PD=2.35657e-06 PS=1.92657e-06 $X=5800 $Y=2410 $dt=1
M14 Q 8 vdd3i! vdd3i! pe3i L=3.00021e-07 W=1.42657e-06 AD=3.433e-13 AS=4.866e-13 PD=1.92657e-06 PS=2.35657e-06 $X=6640 $Y=2410 $dt=1
M15 vdd3i! 8 Q vdd3i! pe3i L=3.00021e-07 W=1.42657e-06 AD=8.562e-13 AS=3.433e-13 PD=4.53657e-06 PS=1.92657e-06 $X=7480 $Y=2410 $dt=1
.ends ON21JI3VX4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND2JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND2JI3VX1 vdd3i! gnd3i! A B Q
*.DEVICECLIMB
** N=8 EP=5 FDC=6
M0 7 A 8 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=2.688e-13 PD=8.1e-07 PS=2.08e-06 $X=820 $Y=990 $dt=0
M1 gnd3i! B 7 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=2.57137e-13 AS=7e-14 PD=1.43669e-06 PS=8.1e-07 $X=1420 $Y=990 $dt=0
M2 Q 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=4.08663e-13 PD=2.74e-06 PS=2.28331e-06 $X=2390 $Y=660 $dt=0
M3 8 A vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=7.276e-13 PD=1.24e-06 PS=4.56e-06 $X=580 $Y=2410 $dt=1
M4 vdd3i! B 8 vdd3i! pe3i L=3e-07 W=7e-07 AD=3.64829e-13 AS=1.89e-13 PD=1.6455e-06 PS=1.24e-06 $X=1420 $Y=2410 $dt=1
M5 Q 8 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=7.34871e-13 PD=3.78e-06 PS=3.3145e-06 $X=2440 $Y=2410 $dt=1
.ends AND2JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA4JI3VX2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA4JI3VX2 vdd3i! gnd3i! Q D C B A
*.DEVICECLIMB
** N=14 EP=7 FDC=16
M0 14 D gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.78e-13 AS=6.098e-13 PD=1.29e-06 PS=3.52e-06 $X=660 $Y=660 $dt=0
M1 13 C 14 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.8245e-13 AS=1.78e-13 PD=1.3e-06 PS=1.29e-06 $X=1410 $Y=660 $dt=0
M2 12 B 13 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.78e-13 AS=1.8245e-13 PD=1.29e-06 PS=1.3e-06 $X=2170 $Y=660 $dt=0
M3 Q A 12 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.293e-13 AS=1.78e-13 PD=1.63e-06 PS=1.29e-06 $X=2920 $Y=660 $dt=0
M4 11 A Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.78e-13 AS=3.293e-13 PD=1.29e-06 PS=1.63e-06 $X=4010 $Y=660 $dt=0
M5 10 B 11 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.8245e-13 AS=1.78e-13 PD=1.3e-06 PS=1.29e-06 $X=4760 $Y=660 $dt=0
M6 9 C 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.78e-13 AS=1.8245e-13 PD=1.29e-06 PS=1.3e-06 $X=5520 $Y=660 $dt=0
M7 gnd3i! D 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=6.098e-13 AS=1.78e-13 PD=3.52e-06 PS=1.29e-06 $X=6270 $Y=660 $dt=0
M8 vdd3i! D Q vdd3i! pe3i L=3.00056e-07 W=9.91066e-07 AD=6.12287e-13 AS=4.22737e-13 PD=2.90357e-06 PS=2.83607e-06 $X=620 $Y=2410 $dt=1
M9 vdd3i! C Q vdd3i! pe3i L=3.00056e-07 W=9.91066e-07 AD=6.12287e-13 AS=2.21137e-13 PD=2.90357e-06 PS=1.45607e-06 $X=1440 $Y=2410 $dt=1
M10 Q B vdd3i! vdd3i! pe3i L=3.00056e-07 W=9.91066e-07 AD=2.21137e-13 AS=6.12287e-13 PD=1.45607e-06 PS=2.90357e-06 $X=2280 $Y=2410 $dt=1
M11 vdd3i! A Q vdd3i! pe3i L=3.00056e-07 W=9.91066e-07 AD=6.12287e-13 AS=2.93137e-13 PD=2.90357e-06 PS=1.60607e-06 $X=2995 $Y=2410 $dt=1
M12 Q A vdd3i! vdd3i! pe3i L=3.00056e-07 W=9.91066e-07 AD=2.93137e-13 AS=6.12287e-13 PD=1.60607e-06 PS=2.90357e-06 $X=3985 $Y=2410 $dt=1
M13 vdd3i! B Q vdd3i! pe3i L=3.00056e-07 W=9.91066e-07 AD=6.12287e-13 AS=2.21137e-13 PD=2.90357e-06 PS=1.45607e-06 $X=4700 $Y=2410 $dt=1
M14 Q C vdd3i! vdd3i! pe3i L=3.00056e-07 W=9.91066e-07 AD=2.21137e-13 AS=6.12287e-13 PD=1.45607e-06 PS=2.90357e-06 $X=5540 $Y=2410 $dt=1
M15 Q D vdd3i! vdd3i! pe3i L=3.00056e-07 W=9.91066e-07 AD=4.22737e-13 AS=6.12287e-13 PD=2.83607e-06 PS=2.90357e-06 $X=6360 $Y=2410 $dt=1
.ends NA4JI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO2I1JI3VX2                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO2I1JI3VX2 vdd3i! gnd3i! AN Q B
*.DEVICECLIMB
** N=9 EP=5 FDC=10
M0 gnd3i! AN 7 gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.3695e-13 AS=4.15012e-13 PD=1.44536e-06 PS=2.72536e-06 $X=595 $Y=660 $dt=0
M1 Q 7 gnd3i! gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.28113e-13 AS=2.3695e-13 PD=1.41536e-06 PS=1.44536e-06 $X=1500 $Y=660 $dt=0
M2 gnd3i! B Q gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.30162e-13 AS=2.28113e-13 PD=1.43036e-06 PS=1.41536e-06 $X=2340 $Y=660 $dt=0
M3 Q B gnd3i! gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.28113e-13 AS=2.30162e-13 PD=1.41536e-06 PS=1.43036e-06 $X=3230 $Y=660 $dt=0
M4 gnd3i! 7 Q gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=4.20212e-13 AS=2.28113e-13 PD=2.75536e-06 PS=1.41536e-06 $X=4070 $Y=660 $dt=0
M5 vdd3i! AN 7 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.998e-13 AS=6.768e-13 PD=2.595e-06 PS=3.78e-06 $X=620 $Y=2410 $dt=1
M6 9 7 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.115e-13 AS=6.998e-13 PD=1.71e-06 PS=2.595e-06 $X=1755 $Y=2410 $dt=1
M7 Q B 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.8775e-13 AS=2.115e-13 PD=1.96e-06 PS=1.71e-06 $X=2355 $Y=2410 $dt=1
M8 8 B Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.115e-13 AS=3.8775e-13 PD=1.71e-06 PS=1.96e-06 $X=3205 $Y=2410 $dt=1
M9 vdd3i! 7 8 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.3642e-12 AS=2.115e-13 PD=5.11e-06 PS=1.71e-06 $X=3805 $Y=2410 $dt=1
.ends NO2I1JI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: EO2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt EO2JI3VX0 vdd3i! gnd3i! B A Q
*.DEVICECLIMB
** N=10 EP=5 FDC=10
M0 8 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.628e-13 PD=9.6e-07 PS=3.52e-06 $X=660 $Y=1130 $dt=0
M1 gnd3i! A 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.0445e-13 AS=1.134e-13 PD=1.34e-06 PS=9.6e-07 $X=1550 $Y=1130 $dt=0
M2 7 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.0445e-13 PD=6.7e-07 PS=1.34e-06 $X=2670 $Y=980 $dt=0
M3 Q A 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.503e-13 AS=5.25e-14 PD=1.15e-06 PS=6.7e-07 $X=3270 $Y=980 $dt=0
M4 gnd3i! 8 Q gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.0464e-12 AS=1.503e-13 PD=4.3e-06 PS=1.15e-06 $X=4200 $Y=1130 $dt=0
M5 10 B vdd3i! vdd3i! pe3i L=3e-07 W=9e-07 AD=1.35e-13 AS=7.175e-13 PD=1.2e-06 PS=4.61e-06 $X=575 $Y=2410 $dt=1
M6 8 A 10 vdd3i! pe3i L=3e-07 W=9e-07 AD=5.38188e-13 AS=1.35e-13 PD=3.13778e-06 PS=1.2e-06 $X=1175 $Y=2410 $dt=1
M7 vdd3i! B 9 vdd3i! pe3i L=3e-07 W=1.3e-06 AD=5.321e-13 AS=5.76588e-13 PD=2.43e-06 PS=3.57778e-06 $X=2795 $Y=2520 $dt=1
M8 9 A vdd3i! vdd3i! pe3i L=3e-07 W=1.3e-06 AD=3.835e-13 AS=5.321e-13 PD=1.89e-06 PS=2.43e-06 $X=3765 $Y=2410 $dt=1
M9 Q 8 9 vdd3i! pe3i L=3e-07 W=1.3e-06 AD=6.565e-13 AS=3.835e-13 PD=3.61e-06 PS=1.89e-06 $X=4655 $Y=2410 $dt=1
.ends EO2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND2JI3VX0                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND2JI3VX0 vdd3i! gnd3i! A B Q
*.DEVICECLIMB
** N=8 EP=5 FDC=6
M0 7 A 8 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=2.688e-13 PD=8.1e-07 PS=2.08e-06 $X=820 $Y=990 $dt=0
M1 gnd3i! B 7 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=3.536e-13 AS=7e-14 PD=2.12571e-06 PS=8.1e-07 $X=1420 $Y=990 $dt=0
M2 Q 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=2.652e-13 PD=1.8e-06 PS=1.59429e-06 $X=2390 $Y=1130 $dt=0
M3 8 A vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=7.276e-13 PD=1.24e-06 PS=4.56e-06 $X=580 $Y=2410 $dt=1
M4 vdd3i! B 8 vdd3i! pe3i L=3e-07 W=7e-07 AD=5.276e-13 AS=1.89e-13 PD=2.48e-06 PS=1.24e-06 $X=1420 $Y=2410 $dt=1
M5 Q 8 vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=3.36e-13 AS=5.276e-13 PD=2.36e-06 PS=2.48e-06 $X=2440 $Y=2410 $dt=1
.ends AND2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AN22JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AN22JI3VX1 vdd3i! gnd3i! B A Q C D
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 10 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=6.098e-13 PD=1.14e-06 PS=3.52e-06 $X=660 $Y=660 $dt=0
M1 Q A 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=1.1125e-13 PD=1.43e-06 PS=1.14e-06 $X=1260 $Y=660 $dt=0
M2 9 C Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=2.403e-13 PD=1.14e-06 PS=1.43e-06 $X=2150 $Y=660 $dt=0
M3 gnd3i! D 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=8.082e-13 AS=1.1125e-13 PD=3.84e-06 PS=1.14e-06 $X=2750 $Y=660 $dt=0
M4 vdd3i! B 11 vdd3i! pe3i L=3.01094e-07 W=1.47213e-06 AD=4.29e-13 AS=6.0945e-13 PD=2.32213e-06 PS=3.77213e-06 $X=660 $Y=2410 $dt=1
M5 11 A vdd3i! vdd3i! pe3i L=3.01094e-07 W=1.47213e-06 AD=4.05825e-13 AS=4.29e-13 PD=2.06213e-06 PS=2.32213e-06 $X=1310 $Y=2410 $dt=1
M6 Q C 11 vdd3i! pe3i L=3.01094e-07 W=1.47213e-06 AD=2.9925e-13 AS=4.05825e-13 PD=1.92213e-06 PS=2.06213e-06 $X=2200 $Y=2410 $dt=1
M7 11 D Q vdd3i! pe3i L=3.01094e-07 W=1.47213e-06 AD=6.252e-13 AS=2.9925e-13 PD=3.77213e-06 PS=1.92213e-06 $X=3100 $Y=2410 $dt=1
.ends AN22JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO2JI3VX2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO2JI3VX2 vdd3i! gnd3i! B A Q
*.DEVICECLIMB
** N=8 EP=5 FDC=8
M0 Q B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=6.842e-13 PD=1.43e-06 PS=3.64e-06 $X=720 $Y=660 $dt=0
M1 gnd3i! A Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=1610 $Y=660 $dt=0
M2 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=2580 $Y=660 $dt=0
M3 gnd3i! B Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=6.098e-13 AS=2.403e-13 PD=3.52e-06 PS=1.43e-06 $X=3470 $Y=660 $dt=0
M4 8 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=1.6898e-12 PD=1.66e-06 PS=5.48e-06 $X=1120 $Y=2410 $dt=1
M5 Q A 8 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=1.7625e-13 PD=1.95e-06 PS=1.66e-06 $X=1670 $Y=2410 $dt=1
M6 7 A Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=3.807e-13 PD=1.66e-06 PS=1.95e-06 $X=2510 $Y=2410 $dt=1
M7 vdd3i! B 7 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.6898e-12 AS=1.7625e-13 PD=5.48e-06 PS=1.66e-06 $X=3060 $Y=2410 $dt=1
.ends NO2JI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AO21JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AO21JI3VX1 vdd3i! gnd3i! B A C Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 9 B gnd3i! gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=5.768e-13 PD=8.1e-07 PS=3.52e-06 $X=660 $Y=990 $dt=0
M1 8 A 9 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=1.708e-13 AS=7e-14 PD=1.17e-06 PS=8.1e-07 $X=1260 $Y=990 $dt=0
M2 gnd3i! C 8 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=3.94626e-13 AS=1.708e-13 PD=1.68386e-06 PS=1.17e-06 $X=2220 $Y=990 $dt=0
M3 Q 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=6.27174e-13 PD=2.74e-06 PS=2.67614e-06 $X=3510 $Y=660 $dt=0
M4 vdd3i! B 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=3.8185e-13 AS=4.08e-13 PD=2.53e-06 PS=2.66e-06 $X=620 $Y=2410 $dt=1
M5 10 A vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=2.295e-13 AS=3.8185e-13 PD=1.39e-06 PS=2.53e-06 $X=1340 $Y=2410 $dt=1
M6 8 C 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.08e-13 AS=2.295e-13 PD=2.66e-06 PS=1.39e-06 $X=2180 $Y=2410 $dt=1
M7 Q 8 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=7.0775e-13 PD=3.78e-06 PS=4.73e-06 $X=3560 $Y=2410 $dt=1
.ends AO21JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA2I1JI3VX2                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA2I1JI3VX2 vdd3i! gnd3i! AN Q B
*.DEVICECLIMB
** N=9 EP=5 FDC=10
M0 gnd3i! AN 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.672e-13 AS=4.272e-13 PD=2.05e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 8 9 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=4.672e-13 PD=1.14e-06 PS=2.05e-06 $X=1780 $Y=660 $dt=0
M2 Q B 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.759e-13 AS=1.1125e-13 PD=1.51e-06 PS=1.14e-06 $X=2380 $Y=660 $dt=0
M3 7 B Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=2.759e-13 PD=1.14e-06 PS=1.51e-06 $X=3350 $Y=660 $dt=0
M4 gnd3i! 9 7 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=7.09e-13 AS=1.1125e-13 PD=3.68e-06 PS=1.14e-06 $X=3950 $Y=660 $dt=0
M5 vdd3i! AN 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=9.9878e-13 AS=6.768e-13 PD=4.57664e-06 PS=3.78e-06 $X=620 $Y=2410 $dt=1
M6 Q 9 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.7e-13 AS=7.08355e-13 PD=1.54e-06 PS=3.24584e-06 $X=1540 $Y=2410 $dt=1
M7 vdd3i! B Q vdd3i! pe3i L=3e-07 W=1e-06 AD=7.08355e-13 AS=2.7e-13 PD=3.24584e-06 PS=1.54e-06 $X=2380 $Y=2410 $dt=1
M8 Q B vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.7e-13 AS=7.08355e-13 PD=1.54e-06 PS=3.24584e-06 $X=3280 $Y=2410 $dt=1
M9 vdd3i! 9 Q vdd3i! pe3i L=3e-07 W=1e-06 AD=7.08355e-13 AS=2.7e-13 PD=3.24584e-06 PS=1.54e-06 $X=4120 $Y=2410 $dt=1
.ends NA2I1JI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA22JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA22JI3VX1 vdd3i! gnd3i! A B C Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 9 A 10 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=2.688e-13 PD=8.1e-07 PS=2.08e-06 $X=620 $Y=990 $dt=0
M1 gnd3i! B 9 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=3.3376e-13 AS=7e-14 PD=1.56028e-06 PS=8.1e-07 $X=1220 $Y=990 $dt=0
M2 8 C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=5.3044e-13 PD=1.14e-06 PS=2.47972e-06 $X=2350 $Y=660 $dt=0
M3 Q 10 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=1.1125e-13 PD=2.74e-06 PS=1.14e-06 $X=2950 $Y=660 $dt=0
M4 10 A vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=7.66562e-13 PD=1.24e-06 PS=3.33273e-06 $X=510 $Y=2410 $dt=1
M5 vdd3i! B 10 vdd3i! pe3i L=3e-07 W=7e-07 AD=7.66562e-13 AS=1.89e-13 PD=3.33273e-06 PS=1.24e-06 $X=1350 $Y=2410 $dt=1
M6 vdd3i! C Q vdd3i! pe3i L=3.00052e-07 W=9.98995e-07 AD=1.09399e-12 AS=2.255e-13 PD=4.75626e-06 PS=1.46899e-06 $X=2190 $Y=2410 $dt=1
M7 Q 10 vdd3i! vdd3i! pe3i L=3.00052e-07 W=9.98995e-07 AD=2.255e-13 AS=1.09399e-12 PD=1.46899e-06 PS=4.75626e-06 $X=3030 $Y=2410 $dt=1
.ends NA22JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MU2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MU2JI3VX0 vdd3i! gnd3i! S IN0 IN1 Q
*.DEVICECLIMB
** N=13 EP=6 FDC=12
M0 gnd3i! S 11 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.5315e-13 AS=2.016e-13 PD=1.165e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 10 IN0 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.5315e-13 PD=6.7e-07 PS=1.165e-06 $X=1550 $Y=965 $dt=0
M2 9 11 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=2150 $Y=965 $dt=0
M3 8 S 9 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=3040 $Y=965 $dt=0
M4 gnd3i! IN1 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.148e-13 AS=5.25e-14 PD=1.88e-06 PS=6.7e-07 $X=3640 $Y=965 $dt=0
M5 Q 9 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=3.148e-13 PD=1.8e-06 PS=1.88e-06 $X=4630 $Y=1130 $dt=0
M6 vdd3i! S 11 vdd3i! pe3i L=3e-07 W=5e-07 AD=1.78281e-13 AS=2.525e-13 PD=1.10156e-06 PS=2.01e-06 $X=645 $Y=2675 $dt=1
M7 13 IN0 vdd3i! vdd3i! pe3i L=3e-07 W=7.8e-07 AD=1.17e-13 AS=2.78119e-13 PD=1.08e-06 PS=1.71844e-06 $X=1575 $Y=2675 $dt=1
M8 9 S 13 vdd3i! pe3i L=3e-07 W=7.8e-07 AD=2.301e-13 AS=1.17e-13 PD=1.37e-06 PS=1.08e-06 $X=2175 $Y=2675 $dt=1
M9 12 11 9 vdd3i! pe3i L=3e-07 W=7.8e-07 AD=1.17e-13 AS=2.301e-13 PD=1.08e-06 PS=1.37e-06 $X=3065 $Y=2675 $dt=1
M10 vdd3i! IN1 12 vdd3i! pe3i L=3e-07 W=7.8e-07 AD=5.0563e-13 AS=1.17e-13 PD=2.58243e-06 PS=1.08e-06 $X=3665 $Y=2675 $dt=1
M11 Q 9 vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=3.535e-13 AS=4.5377e-13 PD=2.41e-06 PS=2.31757e-06 $X=4655 $Y=2410 $dt=1
.ends MU2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OR3JI3VX1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OR3JI3VX1 vdd3i! gnd3i! A B C Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 gnd3i! A 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.482e-13 AS=2.016e-13 PD=2.04e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 8 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.116e-13 AS=2.482e-13 PD=1.78e-06 PS=2.04e-06 $X=1390 $Y=1310 $dt=0
M2 gnd3i! C 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.66689e-13 AS=2.116e-13 PD=1.17398e-06 PS=1.78e-06 $X=2160 $Y=1130 $dt=0
M3 Q 8 gnd3i! gnd3i! ne3i L=3.50112e-07 W=8.98284e-07 AD=4.174e-13 AS=3.56511e-13 PD=2.72828e-06 PS=2.51087e-06 $X=2970 $Y=660 $dt=0
M4 10 A 8 vdd3i! pe3i L=3e-07 W=1e-06 AD=1.375e-13 AS=4.8e-13 PD=1.275e-06 PS=2.96e-06 $X=670 $Y=2720 $dt=1
M5 9 B 10 vdd3i! pe3i L=3e-07 W=1e-06 AD=1.375e-13 AS=1.375e-13 PD=1.275e-06 PS=1.275e-06 $X=1245 $Y=2720 $dt=1
M6 vdd3i! C 9 vdd3i! pe3i L=3e-07 W=1e-06 AD=5.59502e-13 AS=1.375e-13 PD=2.19087e-06 PS=1.275e-06 $X=1820 $Y=2720 $dt=1
M7 Q 8 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=7.88898e-13 PD=3.78e-06 PS=3.08913e-06 $X=3000 $Y=2410 $dt=1
.ends OR3JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ON211JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ON211JI3VX1 vdd3i! gnd3i! B Q A C D
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 Q B 10 gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.27987e-13 AS=4.20337e-13 PD=1.41536e-06 PS=2.75536e-06 $X=620 $Y=660 $dt=0
M1 10 A Q gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.30287e-13 AS=2.27987e-13 PD=1.43036e-06 PS=1.41536e-06 $X=1460 $Y=660 $dt=0
M2 9 C 10 gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=1.21188e-13 AS=2.30287e-13 PD=1.17536e-06 PS=1.43036e-06 $X=2350 $Y=660 $dt=0
M3 gnd3i! D 9 gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=4.20337e-13 AS=1.21188e-13 PD=2.75536e-06 PS=1.17536e-06 $X=2950 $Y=660 $dt=0
M4 11 B vdd3i! vdd3i! pe3i L=3e-07 W=1.38e-06 AD=1.725e-13 AS=9.388e-13 PD=1.63e-06 PS=4.63e-06 $X=695 $Y=2410 $dt=1
M5 Q A 11 vdd3i! pe3i L=3e-07 W=1.38e-06 AD=4.69617e-13 AS=1.725e-13 PD=2.38255e-06 PS=1.63e-06 $X=1245 $Y=2410 $dt=1
M6 vdd3i! C Q vdd3i! pe3i L=3.00049e-07 W=9.66924e-07 AD=4.25413e-13 AS=3.29046e-13 PD=2.34192e-06 PS=1.66938e-06 $X=2210 $Y=2410 $dt=1
M7 Q D vdd3i! vdd3i! pe3i L=3.00049e-07 W=9.66924e-07 AD=4.20162e-13 AS=4.25413e-13 PD=2.80192e-06 PS=2.34192e-06 $X=3000 $Y=2410 $dt=1
.ends ON211JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AN21JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AN21JI3VX1 vdd3i! gnd3i! B A Q C
*.DEVICECLIMB
** N=9 EP=6 FDC=6
M0 8 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=6.47e-13 PD=1.14e-06 PS=3.58e-06 $X=690 $Y=660 $dt=0
M1 Q A 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.28413e-13 AS=1.1125e-13 PD=1.78572e-06 PS=1.14e-06 $X=1290 $Y=660 $dt=0
M2 gnd3i! C Q gnd3i! ne3i L=3.5e-07 W=6.65e-07 AD=6.369e-13 AS=2.45387e-13 PD=3.6e-06 PS=1.33428e-06 $X=2310 $Y=885 $dt=0
M3 vdd3i! B 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.371e-13 AS=6.768e-13 PD=2.03e-06 PS=3.78e-06 $X=620 $Y=2410 $dt=1
M4 9 A vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=4.371e-13 PD=1.95e-06 PS=2.03e-06 $X=1540 $Y=2410 $dt=1
M5 Q C 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.614e-13 AS=3.807e-13 PD=3.9e-06 PS=1.95e-06 $X=2380 $Y=2410 $dt=1
.ends AN21JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INJI3VX0                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INJI3VX0 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=5 EP=4 FDC=2
M0 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=6.248e-13 PD=1.8e-06 PS=3.62e-06 $X=710 $Y=1130 $dt=0
M1 Q A vdd3i! vdd3i! pe3i L=3e-07 W=9.4e-07 AD=4.512e-13 AS=1.0092e-12 PD=2.84e-06 PS=4.76e-06 $X=760 $Y=2410 $dt=1
.ends INJI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO3I1JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO3I1JI3VX1 vdd3i! gnd3i! AN Q B C
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 gnd3i! AN 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.99484e-13 AS=2.016e-13 PD=1.19267e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 Q 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=4.22716e-13 PD=1.43e-06 PS=2.52733e-06 $X=1550 $Y=660 $dt=0
M2 gnd3i! B Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=2440 $Y=660 $dt=0
M3 Q C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=3.494e-13 PD=2.74e-06 PS=1.86e-06 $X=3410 $Y=660 $dt=0
M4 vdd3i! AN 8 vdd3i! pe3i L=3e-07 W=7e-07 AD=4.49443e-13 AS=3.36e-13 PD=1.73175e-06 PS=2.36e-06 $X=620 $Y=2415 $dt=1
M5 10 8 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=9.05307e-13 PD=1.72e-06 PS=3.48825e-06 $X=1770 $Y=2410 $dt=1
M6 9 B 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=2.1855e-13 PD=1.72e-06 PS=1.72e-06 $X=2380 $Y=2410 $dt=1
M7 Q C 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=2.1855e-13 PD=3.78e-06 PS=1.72e-06 $X=2990 $Y=2410 $dt=1
.ends NO3I1JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP25JI3V                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP25JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=12
M0 gnd3i! 5 4 gnd3i! ne3i L=3.5e-07 W=8.8e-07 AD=2.376e-13 AS=4.224e-13 PD=1.42e-06 PS=2.72e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=1510 $Y=660 $dt=0
M2 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=3990 $Y=660 $dt=0
M3 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=6470 $Y=660 $dt=0
M4 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=8950 $Y=660 $dt=0
M5 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=4.312e-13 AS=2.376e-13 PD=2.74e-06 PS=1.42e-06 $X=11430 $Y=660 $dt=0
M6 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.5505e-13 AS=6.312e-13 PD=1.855e-06 PS=3.59e-06 $X=620 $Y=2505 $dt=1
M7 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.5505e-13 AS=3.5505e-13 PD=1.855e-06 PS=1.855e-06 $X=3090 $Y=2505 $dt=1
M8 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.5505e-13 AS=3.5505e-13 PD=1.855e-06 PS=1.855e-06 $X=5560 $Y=2505 $dt=1
M9 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.5505e-13 AS=3.5505e-13 PD=1.855e-06 PS=1.855e-06 $X=8030 $Y=2505 $dt=1
M10 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.84638e-13 AS=3.5505e-13 PD=1.9e-06 PS=1.855e-06 $X=10500 $Y=2505 $dt=1
M11 5 4 vdd3i! vdd3i! pe3i L=3e-07 W=1.315e-06 AD=7.56575e-13 AS=3.84638e-13 PD=3.91e-06 PS=1.9e-06 $X=13015 $Y=2505 $dt=1
.ends DECAP25JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP15JI3V                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP15JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=8
M0 gnd3i! 5 4 gnd3i! ne3i L=3.5e-07 W=8.8e-07 AD=2.42e-13 AS=4.224e-13 PD=1.43e-06 PS=2.72e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.71e-06 W=8.8e-07 AD=2.42e-13 AS=2.42e-13 PD=1.43e-06 PS=1.43e-06 $X=1520 $Y=660 $dt=0
M2 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.71e-06 W=8.8e-07 AD=2.376e-13 AS=2.42e-13 PD=1.42e-06 PS=1.43e-06 $X=3780 $Y=660 $dt=0
M3 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.71e-06 W=8.8e-07 AD=6.046e-13 AS=2.376e-13 PD=3.5e-06 PS=1.42e-06 $X=6030 $Y=660 $dt=0
M4 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.7e-06 W=1.315e-06 AD=3.5505e-13 AS=8.308e-13 PD=1.855e-06 PS=4.37e-06 $X=660 $Y=2505 $dt=1
M5 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.7e-06 W=1.315e-06 AD=3.5505e-13 AS=3.5505e-13 PD=1.855e-06 PS=1.855e-06 $X=2900 $Y=2505 $dt=1
M6 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.7e-06 W=1.315e-06 AD=3.78063e-13 AS=3.5505e-13 PD=1.89e-06 PS=1.855e-06 $X=5140 $Y=2505 $dt=1
M7 5 4 vdd3i! vdd3i! pe3i L=3e-07 W=1.315e-06 AD=7.56575e-13 AS=3.78063e-13 PD=3.91e-06 PS=1.89e-06 $X=7415 $Y=2505 $dt=1
.ends DECAP15JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP7JI3V                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP7JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=4
M0 gnd3i! 5 4 gnd3i! ne3i L=3.5e-07 W=8.8e-07 AD=2.376e-13 AS=4.224e-13 PD=1.42e-06 PS=2.72e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.75e-06 W=8.8e-07 AD=6.046e-13 AS=2.376e-13 PD=3.5e-06 PS=1.42e-06 $X=1510 $Y=660 $dt=0
M2 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.71e-06 W=1.315e-06 AD=3.87925e-13 AS=8.308e-13 PD=1.905e-06 PS=4.37e-06 $X=660 $Y=2505 $dt=1
M3 5 4 vdd3i! vdd3i! pe3i L=3e-07 W=1.315e-06 AD=7.237e-13 AS=3.87925e-13 PD=3.86e-06 PS=1.905e-06 $X=2960 $Y=2505 $dt=1
.ends DECAP7JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP5JI3V                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP5JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=2
M0 gnd3i! 5 4 gnd3i! ne3i L=1.48e-06 W=8.3e-07 AD=5.786e-13 AS=4.568e-13 PD=3.4e-06 PS=2.82e-06 $X=660 $Y=660 $dt=0
M1 5 4 vdd3i! vdd3i! pe3i L=1.46e-06 W=1.36e-06 AD=7.564e-13 AS=8.542e-13 PD=3.9e-06 PS=4.46e-06 $X=660 $Y=2460 $dt=1
.ends DECAP5JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP10JI3V                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP10JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=6
M0 gnd3i! 5 4 gnd3i! ne3i L=3.5e-07 W=8.8e-07 AD=2.376e-13 AS=4.224e-13 PD=1.42e-06 PS=2.72e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.445e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=1510 $Y=660 $dt=0
M2 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.445e-06 W=8.8e-07 AD=6.046e-13 AS=2.376e-13 PD=3.5e-06 PS=1.42e-06 $X=3495 $Y=660 $dt=0
M3 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.425e-06 W=1.315e-06 AD=3.5505e-13 AS=8.308e-13 PD=1.855e-06 PS=4.37e-06 $X=660 $Y=2505 $dt=1
M4 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.425e-06 W=1.315e-06 AD=3.71488e-13 AS=3.5505e-13 PD=1.88e-06 PS=1.855e-06 $X=2625 $Y=2505 $dt=1
M5 5 4 vdd3i! vdd3i! pe3i L=3e-07 W=1.315e-06 AD=7.56575e-13 AS=3.71488e-13 PD=3.91e-06 PS=1.88e-06 $X=4615 $Y=2505 $dt=1
.ends DECAP10JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: aska_dig                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt aska_dig DAC<0> DAC<1> DAC<2> DAC<3> DAC<4> DAC<5> IC_addr<0> IC_addr<1> SPI_CS SPI_Clk
+ SPI_MOSI clk down_switches<0> down_switches<10> down_switches<11> down_switches<12> down_switches<13> down_switches<14> down_switches<15> down_switches<16>
+ down_switches<17> down_switches<18> down_switches<19> down_switches<1> down_switches<20> down_switches<21> down_switches<22> down_switches<23> down_switches<24> down_switches<25>
+ down_switches<26> down_switches<27> down_switches<28> down_switches<29> down_switches<2> down_switches<30> down_switches<31> down_switches<3> down_switches<4> down_switches<5>
+ down_switches<6> down_switches<7> down_switches<8> down_switches<9> enable porborn pulse_active reset_l up_switches<0> up_switches<10>
+ up_switches<11> up_switches<12> up_switches<13> up_switches<14> up_switches<15> up_switches<16> up_switches<17> up_switches<18> up_switches<19> up_switches<1>
+ up_switches<20> up_switches<21> up_switches<22> up_switches<23> up_switches<24> up_switches<25> up_switches<26> up_switches<27> up_switches<28> up_switches<29>
+ up_switches<2> up_switches<30> up_switches<31> up_switches<3> up_switches<4> up_switches<5> up_switches<6> up_switches<7> up_switches<8> up_switches<9>
** N=1434 EP=80 FDC=26952
X8325 1364 1362 80 1155 88 EN2JI3VX0 $T=40320 185920 1 0 $X=39890 $Y=180800
X8326 1364 1362 91 652 701 EN2JI3VX0 $T=45920 185920 1 0 $X=45490 $Y=180800
X8327 1364 1362 498 489 874 EN2JI3VX0 $T=306880 212800 1 180 $X=300850 $Y=212160
X8328 1364 1362 1117 559 1301 565 NO3JI3VX1 $T=347760 24640 1 180 $X=343970 $Y=24000
X8329 1364 1362 480 28 1104 NA2JI3VX2 $T=307440 105280 0 0 $X=307010 $Y=104640
X8330 1364 1362 1096 532 1277 528 NO22JI3VX1 $T=328160 168000 0 180 $X=323250 $Y=162880
X8331 1364 1362 925 607 1141 1365 NO22JI3VX1 $T=397040 141120 1 180 $X=392130 $Y=140480
X8332 1364 1362 533 1111 33 536 DFRRQJI3VX2 $T=342720 212800 0 180 $X=326050 $Y=207680
X8333 1364 1362 1366 DAC<0> BUJI3VX8 $T=50960 33600 1 0 $X=50530 $Y=28480
X8334 1364 1362 1367 DAC<4> BUJI3VX8 $T=67200 33600 1 0 $X=66770 $Y=28480
X8335 1364 1362 152 181 BUJI3VX8 $T=91280 141120 1 0 $X=90850 $Y=136000
X8336 1364 1362 152 180 BUJI3VX8 $T=103600 168000 1 0 $X=103170 $Y=162880
X8337 1364 1362 191 1 BUJI3VX8 $T=126560 203840 0 180 $X=117730 $Y=198720
X8338 1364 1362 191 9 BUJI3VX8 $T=175280 114240 0 0 $X=174850 $Y=113600
X8339 1364 1362 287 DAC<5> BUJI3VX8 $T=176400 24640 1 0 $X=175970 $Y=19520
X8340 1364 1362 191 15 BUJI3VX8 $T=218400 203840 0 0 $X=217970 $Y=203200
X8341 1364 1362 191 19 BUJI3VX8 $T=314720 194880 1 0 $X=314290 $Y=189760
X8342 1364 1362 379 1321 15 456 DFRRQJI3VX4 $T=297360 176960 1 180 $X=279010 $Y=176320
X8343 1364 1362 533 563 33 566 DFRRQJI3VX4 $T=334880 203840 1 0 $X=334450 $Y=198720
X8344 1364 1362 22 914 19 909 DFRRQJI3VX4 $T=379120 185920 1 180 $X=360770 $Y=185280
X8345 1364 1362 22 594 19 606 DFRRQJI3VX4 $T=371840 168000 0 0 $X=371410 $Y=167360
X8346 1364 1362 22 928 19 1139 DFRRQJI3VX4 $T=407680 168000 1 180 $X=389330 $Y=167360
X8347 1364 1362 22 933 19 615 DFRRQJI3VX4 $T=413840 123200 1 180 $X=395490 $Y=122560
X8348 1364 1362 22 1299 19 639 DFRRQJI3VX4 $T=416080 123200 0 180 $X=397730 $Y=118080
X8349 1364 1362 688 723 BUJI3VX1 $T=36960 176960 0 0 $X=36530 $Y=176320
X8350 1364 1362 SPI_Clk 436 BUJI3VX1 $T=120400 96320 0 0 $X=119970 $Y=95680
X8351 1364 1362 clk 555 BUJI3VX1 $T=186480 159040 0 0 $X=186050 $Y=158400
X8352 1364 1362 41 26 BUJI3VX1 $T=207200 87360 1 0 $X=206770 $Y=82240
X8353 1364 1362 350 41 BUJI3VX1 $T=207200 212800 0 0 $X=206770 $Y=212160
X8354 1364 1362 467 44 BUJI3VX1 $T=208320 194880 1 0 $X=207890 $Y=189760
X8355 1364 1362 1041 812 BUJI3VX1 $T=211120 194880 1 0 $X=210690 $Y=189760
X8356 1364 1362 436 688 BUJI3VX1 $T=270480 203840 0 180 $X=267250 $Y=198720
X8357 1364 1362 555 433 BUJI3VX1 $T=339360 185920 0 180 $X=336130 $Y=180800
X8358 1364 1362 462 636 BUJI3VX1 $T=403760 105280 0 0 $X=403330 $Y=104640
X8359 1364 1362 664 45 341 246 NO3I2JI3VX1 $T=209440 185920 1 180 $X=205090 $Y=185280
X8360 1364 1362 14 810 51 1087 NO3I2JI3VX1 $T=220080 176960 0 0 $X=219650 $Y=176320
X8361 1364 1362 197 204 981 183 744 FAJI3VX1 $T=112000 168000 1 0 $X=111570 $Y=162880
X8362 1364 1362 755 744 979 973 187 FAJI3VX1 $T=129360 159040 1 180 $X=114370 $Y=158400
X8363 1364 1362 754 187 223 759 193 FAJI3VX1 $T=133840 150080 0 180 $X=118850 $Y=144960
X8364 1364 1362 976 207 980 757 204 FAJI3VX1 $T=123200 185920 0 0 $X=122770 $Y=185280
X8365 1364 1362 987 208 749 772 199 FAJI3VX1 $T=137760 212800 0 180 $X=122770 $Y=207680
X8366 1364 1362 991 199 978 188 207 FAJI3VX1 $T=141120 203840 0 180 $X=126130 $Y=198720
X8367 1364 1362 235 1196 249 759 244 FAJI3VX1 $T=150640 150080 0 180 $X=135650 $Y=144960
X8368 1364 1362 1202 936 229 973 1196 FAJI3VX1 $T=150640 150080 1 180 $X=135650 $Y=149440
X8369 1364 1362 765 225 217 183 936 FAJI3VX1 $T=151200 168000 0 180 $X=136210 $Y=162880
X8370 1364 1362 219 228 36 757 225 FAJI3VX1 $T=137760 185920 0 0 $X=137330 $Y=185280
X8371 1364 1362 992 767 1200 772 232 FAJI3VX1 $T=140560 212800 0 0 $X=140130 $Y=212160
X8372 1364 1362 1004 232 993 188 228 FAJI3VX1 $T=155680 203840 0 180 $X=140690 $Y=198720
X8373 1364 1362 242 775 771 1368 257 FAJI3VX1 $T=148400 114240 0 0 $X=147970 $Y=113600
X8374 1364 1362 778 193 236 234 274 FAJI3VX1 $T=164640 141120 1 180 $X=149650 $Y=140480
X8375 1364 1362 259 244 771 234 275 FAJI3VX1 $T=166320 150080 1 180 $X=151330 $Y=149440
X8376 1364 1362 784 257 262 253 1015 FAJI3VX1 $T=175840 123200 0 180 $X=160850 $Y=118080
X8377 1364 1362 1306 274 264 258 284 FAJI3VX1 $T=180320 141120 0 180 $X=165330 $Y=136000
X8378 1364 1362 781 275 262 258 289 FAJI3VX1 $T=181440 150080 1 180 $X=166450 $Y=149440
X8379 1364 1362 795 299 800 OR2JI3VX0 $T=183680 194880 0 0 $X=183250 $Y=194240
X8380 1364 1362 360 140 47 OR2JI3VX0 $T=208880 168000 0 0 $X=208450 $Y=167360
X8381 1364 1362 385 1073 1069 OR2JI3VX0 $T=240800 168000 0 0 $X=240370 $Y=167360
X8382 1364 1362 487 140 1270 OR2JI3VX0 $T=303520 168000 1 0 $X=303090 $Y=162880
X8383 1364 1362 384 553 641 OR2JI3VX0 $T=388080 159040 1 0 $X=387650 $Y=153920
X8384 1364 1362 81 1369 78 83 NA3I1JI3VX1 $T=36960 150080 0 0 $X=36530 $Y=149440
X8385 1364 1362 714 1353 956 957 NA3I1JI3VX1 $T=61040 176960 0 0 $X=60610 $Y=176320
X8386 1364 1362 712 482 121 1370 NA3I1JI3VX1 $T=64400 168000 1 0 $X=63970 $Y=162880
X8387 1364 1362 711 712 713 97 NA3I1JI3VX1 $T=68880 159040 1 180 $X=64530 $Y=158400
X8388 1364 1362 536 499 519 557 NA3I1JI3VX1 $T=329280 212800 1 180 $X=324930 $Y=212160
X8389 1364 1362 892 1282 525 888 NA3I1JI3VX1 $T=337680 168000 0 180 $X=333330 $Y=162880
X8390 1364 1362 606 1371 628 1139 NA3I1JI3VX1 $T=386960 168000 1 0 $X=386530 $Y=162880
X8391 1364 1362 615 1372 639 626 NA3I1JI3VX1 $T=395920 114240 1 180 $X=391570 $Y=113600
X8392 1364 1362 636 931 1147 639 NA3I1JI3VX1 $T=401520 114240 1 0 $X=401090 $Y=109120
X8393 1364 1362 152 170 DLY2JI3VX1 $T=77840 212800 0 0 $X=77410 $Y=212160
X8394 1364 1362 70 81 1154 68 NA3JI3VX0 $T=40320 168000 0 180 $X=37090 $Y=162880
X8395 1364 1362 1373 96 704 27 NA3JI3VX0 $T=57120 159040 1 180 $X=53890 $Y=158400
X8396 1364 1362 1374 114 105 113 NA3JI3VX0 $T=58240 150080 0 0 $X=57810 $Y=149440
X8397 1364 1362 70 4 129 132 NA3JI3VX0 $T=67760 185920 0 0 $X=67330 $Y=185280
X8398 1364 1362 132 118 720 122 NA3JI3VX0 $T=75600 194880 0 180 $X=72370 $Y=189760
X8399 1364 1362 982 758 988 227 NA3JI3VX0 $T=133280 123200 1 0 $X=132850 $Y=118080
X8400 1364 1362 222 220 1375 7 NA3JI3VX0 $T=141120 114240 0 0 $X=140690 $Y=113600
X8401 1364 1362 38 774 37 1008 NA3JI3VX0 $T=154560 105280 0 0 $X=154130 $Y=104640
X8402 1364 1362 315 288 317 45 NA3JI3VX0 $T=194320 176960 0 180 $X=191090 $Y=171840
X8403 1364 1362 1033 1031 318 1219 NA3JI3VX0 $T=194320 185920 1 180 $X=191090 $Y=185280
X8404 1364 1362 1032 334 803 1037 NA3JI3VX0 $T=196560 203840 1 0 $X=196130 $Y=198720
X8405 1364 1362 1153 370 834 52 NA3JI3VX0 $T=240800 185920 1 180 $X=237570 $Y=185280
X8406 1364 1362 1376 407 402 405 NA3JI3VX0 $T=250320 159040 0 0 $X=249890 $Y=158400
X8407 1364 1362 45 423 856 858 NA3JI3VX0 $T=271040 185920 1 0 $X=270610 $Y=180800
X8408 1364 1362 78 96 1159 943 ON21JI3VX1 $T=36960 159040 0 180 $X=33170 $Y=153920
X8409 1364 1362 70 1159 1160 703 ON21JI3VX1 $T=38640 159040 1 0 $X=38210 $Y=153920
X8410 1364 1362 1172 117 1302 708 ON21JI3VX1 $T=62720 168000 1 180 $X=58930 $Y=167360
X8411 1364 1362 129 139 1304 4 ON21JI3VX1 $T=72800 185920 0 0 $X=72370 $Y=185280
X8412 1364 1362 292 1377 1215 798 ON21JI3VX1 $T=180880 176960 0 0 $X=180450 $Y=176320
X8413 1364 1362 1378 288 1333 797 ON21JI3VX1 $T=191520 168000 1 180 $X=187730 $Y=167360
X8414 1364 1362 1034 1029 802 318 ON21JI3VX1 $T=194320 185920 1 0 $X=193890 $Y=180800
X8415 1364 1362 47 808 1310 1229 ON21JI3VX1 $T=202720 168000 1 0 $X=202290 $Y=162880
X8416 1364 1362 140 356 1379 1227 ON21JI3VX1 $T=209440 176960 0 180 $X=205650 $Y=171840
X8417 1364 1362 1045 48 358 807 ON21JI3VX1 $T=210560 185920 0 0 $X=210130 $Y=185280
X8418 1364 1362 1055 1335 827 1233 ON21JI3VX1 $T=218960 203840 1 0 $X=218530 $Y=198720
X8419 1364 1362 834 1070 1235 370 ON21JI3VX1 $T=237440 185920 1 180 $X=233650 $Y=185280
X8420 1364 1362 837 1063 1380 1069 ON21JI3VX1 $T=241920 159040 0 0 $X=241490 $Y=158400
X8421 1364 1362 1068 405 1071 840 ON21JI3VX1 $T=249760 168000 0 180 $X=245970 $Y=162880
X8422 1364 1362 404 836 845 1075 ON21JI3VX1 $T=250320 168000 0 0 $X=249890 $Y=167360
X8423 1364 1362 384 848 527 1320 ON21JI3VX1 $T=258160 33600 0 0 $X=257730 $Y=32960
X8424 1364 1362 140 1087 1381 1227 ON21JI3VX1 $T=264880 176960 0 0 $X=264450 $Y=176320
X8425 1364 1362 1382 423 1321 452 ON21JI3VX1 $T=285600 185920 0 180 $X=281810 $Y=180800
X8426 1364 1362 384 866 549 859 ON21JI3VX1 $T=283920 33600 0 0 $X=283490 $Y=32960
X8427 1364 1362 384 470 869 865 ON21JI3VX1 $T=285040 24640 0 0 $X=284610 $Y=24000
X8428 1364 1362 881 1383 500 1273 ON21JI3VX1 $T=317520 168000 1 180 $X=313730 $Y=167360
X8429 1364 1362 384 56 898 1287 ON21JI3VX1 $T=337680 33600 0 0 $X=337250 $Y=32960
X8430 1364 1362 384 1384 908 906 ON21JI3VX1 $T=348880 42560 1 0 $X=348450 $Y=37440
X8431 1364 1362 1121 903 914 60 ON21JI3VX1 $T=360080 185920 1 0 $X=359650 $Y=180800
X8432 1364 1362 384 1349 1126 1348 ON21JI3VX1 $T=371280 33600 1 180 $X=367490 $Y=32960
X8433 1364 1362 384 1135 603 1327 ON21JI3VX1 $T=376880 24640 0 0 $X=376450 $Y=24000
X8434 1364 1362 1371 941 594 610 ON21JI3VX1 $T=384720 168000 0 180 $X=380930 $Y=162880
X8435 1364 1362 1139 1352 1385 631 ON21JI3VX1 $T=390880 159040 1 180 $X=387090 $Y=158400
X8436 1364 1362 627 1365 919 625 ON21JI3VX1 $T=391440 141120 1 180 $X=387650 $Y=140480
X8437 1364 1362 1386 621 1351 615 ON21JI3VX1 $T=388640 114240 0 0 $X=388210 $Y=113600
X8438 1364 1362 628 1352 1146 641 ON21JI3VX1 $T=392000 159040 1 0 $X=391570 $Y=153920
X8439 1364 1362 1372 63 933 1351 ON21JI3VX1 $T=397600 114240 0 0 $X=397170 $Y=113600
X8440 1364 1362 639 63 1299 931 ON21JI3VX1 $T=403760 114240 0 0 $X=403330 $Y=113600
X8441 1364 1362 959 957 714 117 OA21JI3VX1 $T=69440 176960 1 180 $X=64530 $Y=176320
X8442 1364 1362 489 509 520 1106 OA21JI3VX1 $T=316400 212800 0 0 $X=315970 $Y=212160
X8443 1364 1362 152 166 BUJI3VX3 $T=110320 203840 1 0 $X=109890 $Y=198720
X8444 1364 1362 152 169 BUJI3VX3 $T=113680 212800 1 0 $X=113250 $Y=207680
X8445 1364 1362 152 975 BUJI3VX3 $T=119280 212800 1 0 $X=118850 $Y=207680
X8446 1364 1362 152 211 BUJI3VX3 $T=136640 176960 1 0 $X=136210 $Y=171840
X8447 1364 1362 152 213 BUJI3VX3 $T=137200 168000 0 0 $X=136770 $Y=167360
X8448 1364 1362 152 206 BUJI3VX3 $T=137760 185920 1 0 $X=137330 $Y=180800
X8449 1364 1362 152 339 BUJI3VX3 $T=189280 159040 0 0 $X=188850 $Y=158400
X8450 1364 1362 330 up_switches<0> BUJI3VX3 $T=203840 24640 1 0 $X=203410 $Y=19520
X8451 1364 1362 348 up_switches<9> BUJI3VX3 $T=208880 24640 1 0 $X=208450 $Y=19520
X8452 1364 1362 357 up_switches<8> BUJI3VX3 $T=213360 24640 1 0 $X=212930 $Y=19520
X8453 1364 1362 338 up_switches<6> BUJI3VX3 $T=213360 24640 0 0 $X=212930 $Y=24000
X8454 1364 1362 365 up_switches<3> BUJI3VX3 $T=221200 24640 1 180 $X=216850 $Y=24000
X8455 1364 1362 141 up_switches<2> BUJI3VX3 $T=217840 24640 1 0 $X=217410 $Y=19520
X8456 1364 1362 152 822 BUJI3VX3 $T=220640 168000 1 0 $X=220210 $Y=162880
X8457 1364 1362 369 406 BUJI3VX3 $T=220640 194880 1 0 $X=220210 $Y=189760
X8458 1364 1362 152 819 BUJI3VX3 $T=234640 150080 0 180 $X=230290 $Y=144960
X8459 1364 1362 406 467 BUJI3VX3 $T=233520 176960 1 0 $X=233090 $Y=171840
X8460 1364 1362 142 up_switches<1> BUJI3VX3 $T=240800 24640 1 0 $X=240370 $Y=19520
X8461 1364 1362 388 up_switches<4> BUJI3VX3 $T=245840 24640 1 0 $X=245410 $Y=19520
X8462 1364 1362 398 up_switches<10> BUJI3VX3 $T=253120 24640 1 0 $X=252690 $Y=19520
X8463 1364 1362 152 391 BUJI3VX3 $T=255360 123200 0 0 $X=254930 $Y=122560
X8464 1364 1362 342 up_switches<7> BUJI3VX3 $T=258720 24640 1 0 $X=258290 $Y=19520
X8465 1364 1362 422 up_switches<5> BUJI3VX3 $T=264880 24640 1 0 $X=264450 $Y=19520
X8466 1364 1362 439 up_switches<12> BUJI3VX3 $T=271600 24640 1 0 $X=271170 $Y=19520
X8467 1364 1362 283 up_switches<11> BUJI3VX3 $T=277200 24640 1 0 $X=276770 $Y=19520
X8468 1364 1362 354 up_switches<13> BUJI3VX3 $T=282240 24640 1 0 $X=281810 $Y=19520
X8469 1364 1362 692 951 92 90 1161 AN211JI3VX1 $T=45360 168000 0 0 $X=44930 $Y=167360
X8470 1364 1362 105 711 1373 140 116 AN211JI3VX1 $T=64400 159040 1 180 $X=59490 $Y=158400
X8471 1364 1362 1387 272 804 1034 1388 AN211JI3VX1 $T=193200 176960 0 0 $X=192770 $Y=176320
X8472 1364 1362 358 49 341 1057 360 AN211JI3VX1 $T=217280 185920 0 180 $X=212370 $Y=180800
X8473 1364 1362 561 556 1273 562 58 AN211JI3VX1 $T=343280 168000 0 180 $X=338370 $Y=162880
X8474 1364 1362 152 178 BUJI3VX16 $T=110320 203840 0 180 $X=93650 $Y=198720
X8475 1364 1362 777 312 BUJI3VX16 $T=159600 203840 1 0 $X=159170 $Y=198720
X8476 1364 1362 152 320 BUJI3VX16 $T=210000 123200 1 0 $X=209570 $Y=118080
X8477 1364 1362 152 233 BUJI3VX16 $T=239680 132160 0 180 $X=223010 $Y=127040
X8478 1364 1362 71 83 BUJI3VX0 $T=44240 150080 0 0 $X=43810 $Y=149440
X8479 1364 1362 86 950 BUJI3VX0 $T=44240 159040 1 0 $X=43810 $Y=153920
X8480 1364 1362 91 953 BUJI3VX0 $T=54880 194880 1 0 $X=54450 $Y=189760
X8481 1364 1362 654 955 BUJI3VX0 $T=62720 185920 1 0 $X=62290 $Y=180800
X8482 1364 1362 770 1201 BUJI3VX0 $T=151200 114240 1 0 $X=150770 $Y=109120
X8483 1364 1362 776 1355 BUJI3VX0 $T=161840 114240 1 0 $X=161410 $Y=109120
X8484 1364 1362 774 256 BUJI3VX0 $T=162400 96320 1 0 $X=161970 $Y=91200
X8485 1364 1362 243 269 BUJI3VX0 $T=165760 212800 1 0 $X=165330 $Y=207680
X8486 1364 1362 779 1011 BUJI3VX0 $T=190400 105280 0 0 $X=189970 $Y=104640
X8487 1364 1362 44 1041 BUJI3VX0 $T=204960 194880 0 0 $X=204530 $Y=194240
X8488 1364 1362 812 367 BUJI3VX0 $T=207760 194880 0 0 $X=207330 $Y=194240
X8489 1364 1362 815 1313 BUJI3VX0 $T=213920 194880 1 0 $X=213490 $Y=189760
X8490 1364 1362 1313 816 BUJI3VX0 $T=215040 203840 1 0 $X=214610 $Y=198720
X8491 1364 1362 821 815 BUJI3VX0 $T=215600 203840 0 0 $X=215170 $Y=203200
X8492 1364 1362 porborn 821 BUJI3VX0 $T=218400 212800 0 0 $X=217970 $Y=212160
X8493 1364 1362 1072 369 BUJI3VX0 $T=231840 203840 1 0 $X=231410 $Y=198720
X8494 1364 1362 377 52 BUJI3VX0 $T=238000 176960 1 0 $X=237570 $Y=171840
X8495 1364 1362 833 838 BUJI3VX0 $T=241920 203840 0 0 $X=241490 $Y=203200
X8496 1364 1362 843 842 BUJI3VX0 $T=244720 185920 0 0 $X=244290 $Y=185280
X8497 1364 1362 838 1072 BUJI3VX0 $T=244720 212800 1 0 $X=244290 $Y=207680
X8498 1364 1362 SPI_MOSI 1252 BUJI3VX0 $T=260400 212800 0 0 $X=259970 $Y=212160
X8499 1364 1362 852 833 BUJI3VX0 $T=264320 212800 1 0 $X=263890 $Y=207680
X8500 1364 1362 472 479 BUJI3VX0 $T=288960 185920 0 0 $X=288530 $Y=185280
X8501 1364 1362 484 871 BUJI3VX0 $T=295680 194880 1 0 $X=295250 $Y=189760
X8502 1364 1362 874 875 BUJI3VX0 $T=302400 203840 0 0 $X=301970 $Y=203200
X8503 1364 1362 502 520 BUJI3VX0 $T=320880 212800 0 0 $X=320450 $Y=212160
X8504 1364 1362 676 1389 BUJI3VX0 $T=349440 212800 0 0 $X=349010 $Y=212160
X8505 1364 1362 1155 946 80 NA2I1JI3VX1 $T=47600 176960 1 180 $X=43810 $Y=176320
X8506 1364 1362 652 1155 91 NA2I1JI3VX1 $T=50960 176960 1 180 $X=47170 $Y=176320
X8507 1364 1362 100 113 703 NA2I1JI3VX1 $T=57680 150080 1 180 $X=53890 $Y=149440
X8508 1364 1362 703 105 100 NA2I1JI3VX1 $T=54320 159040 1 0 $X=53890 $Y=153920
X8509 1364 1362 1390 710 955 NA2I1JI3VX1 $T=59360 185920 0 0 $X=58930 $Y=185280
X8510 1364 1362 770 999 229 NA2I1JI3VX1 $T=142240 132160 1 0 $X=141810 $Y=127040
X8511 1364 1362 230 1199 999 NA2I1JI3VX1 $T=150080 123200 1 180 $X=146290 $Y=122560
X8512 1364 1362 247 1391 8 NA2I1JI3VX1 $T=160720 132160 0 180 $X=156930 $Y=127040
X8513 1364 1362 779 8 249 NA2I1JI3VX1 $T=162960 123200 1 180 $X=159170 $Y=122560
X8514 1364 1362 1022 791 292 NA2I1JI3VX1 $T=176960 185920 1 0 $X=176530 $Y=180800
X8515 1364 1362 295 318 1035 NA2I1JI3VX1 $T=194880 194880 1 0 $X=194450 $Y=189760
X8516 1364 1362 1035 1037 328 NA2I1JI3VX1 $T=196000 212800 0 0 $X=195570 $Y=212160
X8517 1364 1362 1035 324 295 NA2I1JI3VX1 $T=201600 194880 0 180 $X=197810 $Y=189760
X8518 1364 1362 328 803 1035 NA2I1JI3VX1 $T=199360 203840 1 0 $X=198930 $Y=198720
X8519 1364 1362 340 332 361 NA2I1JI3VX1 $T=204960 176960 0 180 $X=201170 $Y=171840
X8520 1364 1362 14 355 1392 NA2I1JI3VX1 $T=214480 176960 0 180 $X=210690 $Y=171840
X8521 1364 1362 810 666 51 NA2I1JI3VX1 $T=219520 168000 0 0 $X=219090 $Y=167360
X8522 1364 1362 666 487 14 NA2I1JI3VX1 $T=223440 176960 0 180 $X=219650 $Y=171840
X8523 1364 1362 1246 1240 842 NA2I1JI3VX1 $T=250320 194880 0 180 $X=246530 $Y=189760
X8524 1364 1362 446 1393 425 NA2I1JI3VX1 $T=268240 168000 0 180 $X=264450 $Y=162880
X8525 1364 1362 857 438 435 NA2I1JI3VX1 $T=272720 168000 1 180 $X=268930 $Y=167360
X8526 1364 1362 456 435 459 NA2I1JI3VX1 $T=276640 168000 1 180 $X=272850 $Y=167360
X8527 1364 1362 861 425 447 NA2I1JI3VX1 $T=276640 176960 1 180 $X=272850 $Y=176320
X8528 1364 1362 554 518 534 NA2I1JI3VX1 $T=322560 176960 0 180 $X=318770 $Y=171840
X8529 1364 1362 534 529 554 NA2I1JI3VX1 $T=328160 176960 1 0 $X=327730 $Y=171840
X8530 1364 1362 545 900 544 NA2I1JI3VX1 $T=334320 176960 0 0 $X=333890 $Y=176320
X8531 1364 1362 649 944 DLY1JI3VX1 $T=28560 141120 1 0 $X=28130 $Y=136000
X8532 1364 1362 64 687 DLY1JI3VX1 $T=29680 114240 0 0 $X=29250 $Y=113600
X8533 1364 1362 650 686 DLY1JI3VX1 $T=29680 123200 1 0 $X=29250 $Y=118080
X8534 1364 1362 76 689 DLY1JI3VX1 $T=34160 141120 1 0 $X=33730 $Y=136000
X8535 1364 1362 77 690 DLY1JI3VX1 $T=34160 141120 0 0 $X=33730 $Y=140480
X8536 1364 1362 106 1162 DLY1JI3VX1 $T=44240 33600 0 0 $X=43810 $Y=32960
X8537 1364 1362 947 1164 DLY1JI3VX1 $T=47040 123200 0 0 $X=46610 $Y=122560
X8538 1364 1362 651 1166 DLY1JI3VX1 $T=49840 33600 0 0 $X=49410 $Y=32960
X8539 1364 1362 104 1170 DLY1JI3VX1 $T=56000 33600 0 0 $X=55570 $Y=32960
X8540 1364 1362 965 1173 DLY1JI3VX1 $T=61600 33600 0 0 $X=61170 $Y=32960
X8541 1364 1362 1176 961 DLY1JI3VX1 $T=65520 150080 0 0 $X=65090 $Y=149440
X8542 1364 1362 655 1175 DLY1JI3VX1 $T=67200 33600 0 0 $X=66770 $Y=32960
X8543 1364 1362 962 964 DLY1JI3VX1 $T=69440 69440 1 0 $X=69010 $Y=64320
X8544 1364 1362 715 1177 DLY1JI3VX1 $T=72240 141120 0 0 $X=71810 $Y=140480
X8545 1364 1362 138 722 DLY1JI3VX1 $T=72800 33600 0 0 $X=72370 $Y=32960
X8546 1364 1362 656 1179 DLY1JI3VX1 $T=78400 33600 0 0 $X=77970 $Y=32960
X8547 1364 1362 1181 150 DLY1JI3VX1 $T=84560 185920 0 0 $X=84130 $Y=185280
X8548 1364 1362 657 735 DLY1JI3VX1 $T=85120 87360 1 0 $X=84690 $Y=82240
X8549 1364 1362 146 729 DLY1JI3VX1 $T=85120 203840 1 0 $X=84690 $Y=198720
X8550 1364 1362 738 155 DLY1JI3VX1 $T=87360 168000 1 0 $X=86930 $Y=162880
X8551 1364 1362 728 156 DLY1JI3VX1 $T=87360 168000 0 0 $X=86930 $Y=167360
X8552 1364 1362 658 1151 DLY1JI3VX1 $T=89040 150080 1 0 $X=88610 $Y=144960
X8553 1364 1362 731 1180 DLY1JI3VX1 $T=95200 203840 1 180 $X=89170 $Y=203200
X8554 1364 1362 168 1184 DLY1JI3VX1 $T=103040 203840 0 0 $X=102610 $Y=203200
X8555 1364 1362 1182 970 DLY1JI3VX1 $T=103600 69440 0 0 $X=103170 $Y=68800
X8556 1364 1362 1185 972 DLY1JI3VX1 $T=108640 159040 0 0 $X=108210 $Y=158400
X8557 1364 1362 179 974 DLY1JI3VX1 $T=113680 150080 1 0 $X=113250 $Y=144960
X8558 1364 1362 739 745 DLY1JI3VX1 $T=113680 168000 0 0 $X=113250 $Y=167360
X8559 1364 1362 742 748 DLY1JI3VX1 $T=117040 33600 1 0 $X=116610 $Y=28480
X8560 1364 1362 740 985 DLY1JI3VX1 $T=129360 42560 1 0 $X=128930 $Y=37440
X8561 1364 1362 1187 986 DLY1JI3VX1 $T=132160 185920 1 0 $X=131730 $Y=180800
X8562 1364 1362 971 1192 DLY1JI3VX1 $T=134960 42560 1 0 $X=134530 $Y=37440
X8563 1364 1362 1186 990 DLY1JI3VX1 $T=134960 132160 0 0 $X=134530 $Y=131520
X8564 1364 1362 751 762 DLY1JI3VX1 $T=136080 69440 0 0 $X=135650 $Y=68800
X8565 1364 1362 741 995 DLY1JI3VX1 $T=140560 42560 1 0 $X=140130 $Y=37440
X8566 1364 1362 661 1198 DLY1JI3VX1 $T=140560 132160 0 0 $X=140130 $Y=131520
X8567 1364 1362 753 1203 DLY1JI3VX1 $T=146160 42560 1 0 $X=145730 $Y=37440
X8568 1364 1362 998 1003 DLY1JI3VX1 $T=146160 60480 1 0 $X=145730 $Y=55360
X8569 1364 1362 1354 5 DLY1JI3VX1 $T=146160 132160 0 0 $X=145730 $Y=131520
X8570 1364 1362 996 1005 DLY1JI3VX1 $T=151760 60480 1 0 $X=151330 $Y=55360
X8571 1364 1362 764 1205 DLY1JI3VX1 $T=152880 42560 1 0 $X=152450 $Y=37440
X8572 1364 1362 1009 1208 DLY1JI3VX1 $T=157360 60480 1 0 $X=156930 $Y=55360
X8573 1364 1362 1012 1209 DLY1JI3VX1 $T=158480 42560 1 0 $X=158050 $Y=37440
X8574 1364 1362 1016 1018 DLY1JI3VX1 $T=167440 114240 1 0 $X=167010 $Y=109120
X8575 1364 1362 1023 1210 DLY1JI3VX1 $T=169120 33600 0 0 $X=168690 $Y=32960
X8576 1364 1362 1211 1212 DLY1JI3VX1 $T=174720 33600 0 0 $X=174290 $Y=32960
X8577 1364 1362 1020 1309 DLY1JI3VX1 $T=174720 132160 1 0 $X=174290 $Y=127040
X8578 1364 1362 307 1214 DLY1JI3VX1 $T=177520 96320 0 0 $X=177090 $Y=95680
X8579 1364 1362 787 1216 DLY1JI3VX1 $T=179200 42560 1 0 $X=178770 $Y=37440
X8580 1364 1362 1048 1218 DLY1JI3VX1 $T=186480 141120 1 0 $X=186050 $Y=136000
X8581 1364 1362 1036 1220 DLY1JI3VX1 $T=187600 42560 1 0 $X=187170 $Y=37440
X8582 1364 1362 663 1222 DLY1JI3VX1 $T=190960 105280 1 0 $X=190530 $Y=100160
X8583 1364 1362 316 1223 DLY1JI3VX1 $T=192080 33600 0 0 $X=191650 $Y=32960
X8584 1364 1362 1049 1224 DLY1JI3VX1 $T=192080 132160 0 0 $X=191650 $Y=131520
X8585 1364 1362 1030 1225 DLY1JI3VX1 $T=193200 105280 0 0 $X=192770 $Y=104640
X8586 1364 1362 327 336 DLY1JI3VX1 $T=197680 123200 1 0 $X=197250 $Y=118080
X8587 1364 1362 1217 1039 DLY1JI3VX1 $T=197680 132160 0 0 $X=197250 $Y=131520
X8588 1364 1362 SPI_CS 777 DLY1JI3VX1 $T=201600 212800 0 0 $X=201170 $Y=212160
X8589 1364 1362 665 359 DLY1JI3VX1 $T=210000 42560 0 0 $X=209570 $Y=41920
X8590 1364 1362 818 825 DLY1JI3VX1 $T=215600 51520 0 0 $X=215170 $Y=50880
X8591 1364 1362 1064 16 DLY1JI3VX1 $T=217840 42560 1 0 $X=217410 $Y=37440
X8592 1364 1362 1043 1311 DLY1JI3VX1 $T=217840 60480 1 0 $X=217410 $Y=55360
X8593 1364 1362 1236 1237 DLY1JI3VX1 $T=231840 33600 0 0 $X=231410 $Y=32960
X8594 1364 1362 380 1238 DLY1JI3VX1 $T=231840 42560 0 0 $X=231410 $Y=41920
X8595 1364 1362 1312 1062 DLY1JI3VX1 $T=234080 168000 1 0 $X=233650 $Y=162880
X8596 1364 1362 1243 1314 DLY1JI3VX1 $T=235200 168000 0 0 $X=234770 $Y=167360
X8597 1364 1362 1157 667 DLY1JI3VX1 $T=236320 150080 1 0 $X=235890 $Y=144960
X8598 1364 1362 814 387 DLY1JI3VX1 $T=238000 141120 1 0 $X=237570 $Y=136000
X8599 1364 1362 835 1242 DLY1JI3VX1 $T=244160 33600 0 0 $X=243730 $Y=32960
X8600 1364 1362 396 1074 DLY1JI3VX1 $T=245280 141120 1 0 $X=244850 $Y=136000
X8601 1364 1362 1067 1245 DLY1JI3VX1 $T=246960 33600 1 0 $X=246530 $Y=28480
X8602 1364 1362 1254 1079 DLY1JI3VX1 $T=253120 78400 0 0 $X=252690 $Y=77760
X8603 1364 1362 1077 1249 DLY1JI3VX1 $T=254240 42560 0 0 $X=253810 $Y=41920
X8604 1364 1362 420 1081 DLY1JI3VX1 $T=255360 159040 0 0 $X=254930 $Y=158400
X8605 1364 1362 430 1253 DLY1JI3VX1 $T=260960 42560 0 0 $X=260530 $Y=41920
X8606 1364 1362 668 1257 DLY1JI3VX1 $T=265440 150080 1 0 $X=265010 $Y=144960
X8607 1364 1362 442 1258 DLY1JI3VX1 $T=266560 42560 0 0 $X=266130 $Y=41920
X8608 1364 1362 1088 1090 DLY1JI3VX1 $T=270480 168000 1 0 $X=270050 $Y=162880
X8609 1364 1362 1247 1091 DLY1JI3VX1 $T=272160 132160 0 0 $X=271730 $Y=131520
X8610 1364 1362 669 1261 DLY1JI3VX1 $T=273840 42560 0 0 $X=273410 $Y=41920
X8611 1364 1362 1259 1262 DLY1JI3VX1 $T=277760 150080 0 0 $X=277330 $Y=149440
X8612 1364 1362 670 1094 DLY1JI3VX1 $T=283920 69440 0 0 $X=283490 $Y=68800
X8613 1364 1362 476 868 DLY1JI3VX1 $T=286160 168000 0 0 $X=285730 $Y=167360
X8614 1364 1362 473 18 DLY1JI3VX1 $T=288400 114240 0 0 $X=287970 $Y=113600
X8615 1364 1362 1095 1266 DLY1JI3VX1 $T=289520 42560 0 0 $X=289090 $Y=41920
X8616 1364 1362 867 1097 DLY1JI3VX1 $T=289520 69440 0 0 $X=289090 $Y=68800
X8617 1364 1362 870 1267 DLY1JI3VX1 $T=293440 159040 1 0 $X=293010 $Y=153920
X8618 1364 1362 1268 1269 DLY1JI3VX1 $T=297920 42560 0 0 $X=297490 $Y=41920
X8619 1364 1362 671 1271 DLY1JI3VX1 $T=303520 42560 0 0 $X=303090 $Y=41920
X8620 1364 1362 490 495 DLY1JI3VX1 $T=303520 159040 1 0 $X=303090 $Y=153920
X8621 1364 1362 494 1272 DLY1JI3VX1 $T=304640 33600 0 0 $X=304210 $Y=32960
X8622 1364 1362 672 1274 DLY1JI3VX1 $T=309120 42560 0 0 $X=308690 $Y=41920
X8623 1364 1362 1285 1275 DLY1JI3VX1 $T=309680 159040 0 0 $X=309250 $Y=158400
X8624 1364 1362 673 1276 DLY1JI3VX1 $T=315280 42560 0 0 $X=314850 $Y=41920
X8625 1364 1362 521 1323 DLY1JI3VX1 $T=316400 159040 1 0 $X=315970 $Y=153920
X8626 1364 1362 674 1278 DLY1JI3VX1 $T=320880 42560 0 0 $X=320450 $Y=41920
X8627 1364 1362 1103 539 DLY1JI3VX1 $T=327040 42560 1 0 $X=326610 $Y=37440
X8628 1364 1362 1280 540 DLY1JI3VX1 $T=327040 60480 0 0 $X=326610 $Y=59840
X8629 1364 1362 589 1283 DLY1JI3VX1 $T=336000 42560 1 180 $X=329970 $Y=41920
X8630 1364 1362 1114 1288 DLY1JI3VX1 $T=336000 42560 0 0 $X=335570 $Y=41920
X8631 1364 1362 893 1324 DLY1JI3VX1 $T=337680 141120 0 0 $X=337250 $Y=140480
X8632 1364 1362 939 1289 DLY1JI3VX1 $T=347760 176960 0 180 $X=341730 $Y=171840
X8633 1364 1362 675 569 DLY1JI3VX1 $T=342720 51520 0 0 $X=342290 $Y=50880
X8634 1364 1362 1113 1118 DLY1JI3VX1 $T=352240 60480 0 180 $X=346210 $Y=55360
X8635 1364 1362 940 564 DLY1JI3VX1 $T=352240 141120 1 180 $X=346210 $Y=140480
X8636 1364 1362 677 1125 DLY1JI3VX1 $T=360080 150080 1 0 $X=359650 $Y=144960
X8637 1364 1362 1295 1129 DLY1JI3VX1 $T=364560 168000 0 0 $X=364130 $Y=167360
X8638 1364 1362 679 1130 DLY1JI3VX1 $T=365680 150080 1 0 $X=365250 $Y=144960
X8639 1364 1362 1134 916 DLY1JI3VX1 $T=371840 33600 0 0 $X=371410 $Y=32960
X8640 1364 1362 895 1132 DLY1JI3VX1 $T=379120 141120 0 180 $X=373090 $Y=136000
X8641 1364 1362 915 596 DLY1JI3VX1 $T=373520 159040 0 0 $X=373090 $Y=158400
X8642 1364 1362 1133 1296 DLY1JI3VX1 $T=374080 33600 1 0 $X=373650 $Y=28480
X8643 1364 1362 894 599 DLY1JI3VX1 $T=374080 132160 0 0 $X=373650 $Y=131520
X8644 1364 1362 680 605 DLY1JI3VX1 $T=375200 185920 1 0 $X=374770 $Y=180800
X8645 1364 1362 1144 62 DLY1JI3VX1 $T=379680 33600 0 0 $X=379250 $Y=32960
X8646 1364 1362 923 1328 DLY1JI3VX1 $T=385840 24640 1 0 $X=385410 $Y=19520
X8647 1364 1362 922 1298 DLY1JI3VX1 $T=388640 33600 1 0 $X=388210 $Y=28480
X8648 1364 1362 632 1145 DLY1JI3VX1 $T=389760 78400 1 0 $X=389330 $Y=73280
X8649 1364 1362 644 645 DLY1JI3VX1 $T=407680 33600 0 0 $X=407250 $Y=32960
X8650 1364 1362 683 646 DLY1JI3VX1 $T=413280 42560 0 0 $X=412850 $Y=41920
X8651 1364 1362 934 647 DLY1JI3VX1 $T=413280 51520 1 0 $X=412850 $Y=46400
X8652 1364 1362 684 648 DLY1JI3VX1 $T=413280 51520 0 0 $X=412850 $Y=50880
X8653 1364 1362 142 357 306 330 348 OR4JI3VX1 $T=184240 24640 0 0 $X=183810 $Y=24000
X8654 1364 1362 422 388 319 398 283 OR4JI3VX1 $T=199920 24640 0 180 $X=193330 $Y=19520
X8655 1364 1362 342 338 809 439 354 OR4JI3VX1 $T=206080 24640 0 0 $X=205650 $Y=24000
X8656 1364 1362 1126 579 1301 908 898 OR4JI3VX1 $T=366800 24640 1 180 $X=360210 $Y=24000
X8657 1364 1362 72 685 1 68 DFRRQJI3VX1 $T=21280 176960 1 0 $X=20850 $Y=171840
X8658 1364 1362 72 65 1 78 DFRRQJI3VX1 $T=21840 159040 0 0 $X=21410 $Y=158400
X8659 1364 1362 72 66 1 75 DFRRQJI3VX1 $T=21840 185920 1 0 $X=21410 $Y=180800
X8660 1364 1362 72 942 1 71 DFRRQJI3VX1 $T=22400 150080 1 0 $X=21970 $Y=144960
X8661 1364 1362 72 67 1 80 DFRRQJI3VX1 $T=22960 194880 1 0 $X=22530 $Y=189760
X8662 1364 1362 72 73 1 64 DFRRQJI3VX1 $T=39200 105280 0 180 $X=23650 $Y=100160
X8663 1364 1362 72 82 1 649 DFRRQJI3VX1 $T=39760 105280 1 180 $X=24210 $Y=104640
X8664 1364 1362 72 110 1 650 DFRRQJI3VX1 $T=39760 114240 0 180 $X=24210 $Y=109120
X8665 1364 1362 72 687 1 691 DFRRQJI3VX1 $T=24640 123200 0 0 $X=24210 $Y=122560
X8666 1364 1362 72 686 1 693 DFRRQJI3VX1 $T=24640 132160 1 0 $X=24210 $Y=127040
X8667 1364 1362 72 944 1 692 DFRRQJI3VX1 $T=24640 132160 0 0 $X=24210 $Y=131520
X8668 1364 1362 72 950 1 703 DFRRQJI3VX1 $T=39200 150080 1 0 $X=38770 $Y=144960
X8669 1364 1362 72 112 1 76 DFRRQJI3VX1 $T=54880 114240 1 180 $X=39330 $Y=113600
X8670 1364 1362 72 689 1 697 DFRRQJI3VX1 $T=39760 141120 1 0 $X=39330 $Y=136000
X8671 1364 1362 72 690 1 699 DFRRQJI3VX1 $T=39760 141120 0 0 $X=39330 $Y=140480
X8672 1364 1362 72 89 1 91 DFRRQJI3VX1 $T=39760 194880 1 0 $X=39330 $Y=189760
X8673 1364 1362 72 99 1 77 DFRRQJI3VX1 $T=56000 123200 0 180 $X=40450 $Y=118080
X8674 1364 1362 72 95 1 947 DFRRQJI3VX1 $T=57120 132160 0 180 $X=41570 $Y=127040
X8675 1364 1362 72 1164 1 1165 DFRRQJI3VX1 $T=42000 132160 0 0 $X=41570 $Y=131520
X8676 1364 1362 98 1162 1 727 DFRRQJI3VX1 $T=44800 42560 1 0 $X=44370 $Y=37440
X8677 1364 1362 98 1166 1 709 DFRRQJI3VX1 $T=44800 42560 0 0 $X=44370 $Y=41920
X8678 1364 1362 98 84 1 106 DFRRQJI3VX1 $T=44800 51520 1 0 $X=44370 $Y=46400
X8679 1364 1362 98 109 1 651 DFRRQJI3VX1 $T=44800 51520 0 0 $X=44370 $Y=50880
X8680 1364 1362 98 694 1 655 DFRRQJI3VX1 $T=45360 60480 1 0 $X=44930 $Y=55360
X8681 1364 1362 98 695 1 104 DFRRQJI3VX1 $T=45920 69440 1 0 $X=45490 $Y=64320
X8682 1364 1362 72 1168 1 700 DFRRQJI3VX1 $T=62720 194880 1 180 $X=47170 $Y=194240
X8683 1364 1362 72 3 1 654 DFRRQJI3VX1 $T=50960 203840 1 0 $X=50530 $Y=198720
X8684 1364 1362 72 107 1 715 DFRRQJI3VX1 $T=57120 141120 1 0 $X=56690 $Y=136000
X8685 1364 1362 72 1177 1 706 DFRRQJI3VX1 $T=72240 141120 1 180 $X=56690 $Y=140480
X8686 1364 1362 72 961 1 120 DFRRQJI3VX1 $T=72240 150080 0 180 $X=56690 $Y=144960
X8687 1364 1362 72 119 1 122 DFRRQJI3VX1 $T=58240 203840 0 0 $X=57810 $Y=203200
X8688 1364 1362 98 1175 1 721 DFRRQJI3VX1 $T=62160 51520 1 0 $X=61730 $Y=46400
X8689 1364 1362 98 108 1 965 DFRRQJI3VX1 $T=62160 60480 1 0 $X=61730 $Y=55360
X8690 1364 1362 98 1170 1 143 DFRRQJI3VX1 $T=62720 42560 1 0 $X=62290 $Y=37440
X8691 1364 1362 98 1173 1 724 DFRRQJI3VX1 $T=62720 42560 0 0 $X=62290 $Y=41920
X8692 1364 1362 98 958 1 138 DFRRQJI3VX1 $T=63280 60480 0 0 $X=62850 $Y=59840
X8693 1364 1362 98 29 1 656 DFRRQJI3VX1 $T=63840 51520 0 0 $X=63410 $Y=50880
X8694 1364 1362 72 716 1 728 DFRRQJI3VX1 $T=72240 168000 1 0 $X=71810 $Y=162880
X8695 1364 1362 72 156 1 1394 DFRRQJI3VX1 $T=87360 168000 1 180 $X=71810 $Y=167360
X8696 1364 1362 72 935 1 1176 DFRRQJI3VX1 $T=89040 141120 0 180 $X=73490 $Y=136000
X8697 1364 1362 72 1151 1 100 DFRRQJI3VX1 $T=89040 150080 0 180 $X=73490 $Y=144960
X8698 1364 1362 72 1304 1 720 DFRRQJI3VX1 $T=89600 203840 1 180 $X=74050 $Y=203200
X8699 1364 1362 72 150 1 135 DFRRQJI3VX1 $T=90160 185920 0 180 $X=74610 $Y=180800
X8700 1364 1362 72 184 1 731 DFRRQJI3VX1 $T=75040 212800 1 0 $X=74610 $Y=207680
X8701 1364 1362 72 151 1 1181 DFRRQJI3VX1 $T=75600 176960 1 0 $X=75170 $Y=171840
X8702 1364 1362 72 155 1 133 DFRRQJI3VX1 $T=90720 176960 1 180 $X=75170 $Y=176320
X8703 1364 1362 72 967 1 132 DFRRQJI3VX1 $T=90720 194880 1 180 $X=75170 $Y=194240
X8704 1364 1362 98 144 1 962 DFRRQJI3VX1 $T=78400 60480 0 0 $X=77970 $Y=59840
X8705 1364 1362 98 1179 1 153 DFRRQJI3VX1 $T=78960 51520 1 0 $X=78530 $Y=46400
X8706 1364 1362 98 722 1 733 DFRRQJI3VX1 $T=78960 51520 0 0 $X=78530 $Y=50880
X8707 1364 1362 98 964 1 157 DFRRQJI3VX1 $T=78960 60480 1 0 $X=78530 $Y=55360
X8708 1364 1362 98 136 1 657 DFRRQJI3VX1 $T=100240 78400 1 180 $X=84690 $Y=77760
X8709 1364 1362 98 1183 1 658 DFRRQJI3VX1 $T=100240 141120 1 180 $X=84690 $Y=140480
X8710 1364 1362 72 161 1 146 DFRRQJI3VX1 $T=100240 194880 0 180 $X=84690 $Y=189760
X8711 1364 1362 72 1180 1 215 DFRRQJI3VX1 $T=100240 212800 1 180 $X=84690 $Y=212160
X8712 1364 1362 165 748 1 163 DFRRQJI3VX1 $T=98560 42560 1 0 $X=98130 $Y=37440
X8713 1364 1362 165 1192 1 167 DFRRQJI3VX1 $T=98560 42560 0 0 $X=98130 $Y=41920
X8714 1364 1362 98 154 1 742 DFRRQJI3VX1 $T=98560 51520 1 0 $X=98130 $Y=46400
X8715 1364 1362 98 970 1 164 DFRRQJI3VX1 $T=98560 51520 0 0 $X=98130 $Y=50880
X8716 1364 1362 98 969 1 971 DFRRQJI3VX1 $T=98560 60480 1 0 $X=98130 $Y=55360
X8717 1364 1362 98 718 1 1182 DFRRQJI3VX1 $T=98560 60480 0 0 $X=98130 $Y=59840
X8718 1364 1362 72 137 1 739 DFRRQJI3VX1 $T=98560 150080 1 0 $X=98130 $Y=144960
X8719 1364 1362 72 159 1 738 DFRRQJI3VX1 $T=98560 168000 0 0 $X=98130 $Y=167360
X8720 1364 1362 166 162 1 168 DFRRQJI3VX1 $T=98560 194880 0 0 $X=98130 $Y=194240
X8721 1364 1362 169 1184 1 772 DFRRQJI3VX1 $T=98560 212800 1 0 $X=98130 $Y=207680
X8722 1364 1362 170 1197 1 35 DFRRQJI3VX1 $T=100240 212800 0 0 $X=99810 $Y=212160
X8723 1364 1362 98 186 1 1185 DFRRQJI3VX1 $T=102480 123200 1 0 $X=102050 $Y=118080
X8724 1364 1362 98 1188 1 179 DFRRQJI3VX1 $T=103040 132160 0 0 $X=102610 $Y=131520
X8725 1364 1362 178 972 15 973 DFRRQJI3VX1 $T=103600 150080 0 0 $X=103170 $Y=149440
X8726 1364 1362 180 719 1 1187 DFRRQJI3VX1 $T=104160 176960 1 0 $X=103730 $Y=171840
X8727 1364 1362 181 974 1 759 DFRRQJI3VX1 $T=104720 141120 1 0 $X=104290 $Y=136000
X8728 1364 1362 72 745 1 183 DFRRQJI3VX1 $T=104720 176960 0 0 $X=104290 $Y=176320
X8729 1364 1362 975 195 1 749 DFRRQJI3VX1 $T=108640 203840 0 0 $X=108210 $Y=203200
X8730 1364 1362 72 729 1 188 DFRRQJI3VX1 $T=109760 194880 1 0 $X=109330 $Y=189760
X8731 1364 1362 165 735 1 174 DFRRQJI3VX1 $T=128800 51520 1 180 $X=113250 $Y=50880
X8732 1364 1362 165 202 1 741 DFRRQJI3VX1 $T=128800 60480 0 180 $X=113250 $Y=55360
X8733 1364 1362 165 171 1 751 DFRRQJI3VX1 $T=113680 60480 0 0 $X=113250 $Y=59840
X8734 1364 1362 72 660 1 978 DFRRQJI3VX1 $T=113680 194880 0 0 $X=113250 $Y=194240
X8735 1364 1362 165 995 1 192 DFRRQJI3VX1 $T=114240 42560 1 0 $X=113810 $Y=37440
X8736 1364 1362 165 203 1 753 DFRRQJI3VX1 $T=114240 42560 0 0 $X=113810 $Y=41920
X8737 1364 1362 165 1189 1 740 DFRRQJI3VX1 $T=129360 51520 0 180 $X=113810 $Y=46400
X8738 1364 1362 165 985 1 752 DFRRQJI3VX1 $T=114800 33600 0 0 $X=114370 $Y=32960
X8739 1364 1362 98 182 1 1354 DFRRQJI3VX1 $T=118160 114240 0 0 $X=117730 $Y=113600
X8740 1364 1362 98 750 1 1186 DFRRQJI3VX1 $T=133280 123200 0 180 $X=117730 $Y=118080
X8741 1364 1362 98 200 1 661 DFRRQJI3VX1 $T=119840 132160 0 0 $X=119410 $Y=131520
X8742 1364 1362 98 189 1 223 DFRRQJI3VX1 $T=119840 141120 1 0 $X=119410 $Y=136000
X8743 1364 1362 98 190 15 979 DFRRQJI3VX1 $T=119840 150080 0 0 $X=119410 $Y=149440
X8744 1364 1362 206 986 1 757 DFRRQJI3VX1 $T=119840 176960 0 0 $X=119410 $Y=176320
X8745 1364 1362 211 194 1 980 DFRRQJI3VX1 $T=121520 176960 1 0 $X=121090 $Y=171840
X8746 1364 1362 213 1191 1 981 DFRRQJI3VX1 $T=122080 168000 0 0 $X=121650 $Y=167360
X8747 1364 1362 98 990 1 258 DFRRQJI3VX1 $T=123200 132160 1 0 $X=122770 $Y=127040
X8748 1364 1362 165 220 9 198 DFRRQJI3VX1 $T=145600 105280 0 180 $X=130050 $Y=100160
X8749 1364 1362 165 762 9 226 DFRRQJI3VX1 $T=131040 51520 1 0 $X=130610 $Y=46400
X8750 1364 1362 165 1003 9 205 DFRRQJI3VX1 $T=146160 51520 1 180 $X=130610 $Y=50880
X8751 1364 1362 165 1005 9 214 DFRRQJI3VX1 $T=146160 60480 0 180 $X=130610 $Y=55360
X8752 1364 1362 165 209 9 998 DFRRQJI3VX1 $T=131040 60480 0 0 $X=130610 $Y=59840
X8753 1364 1362 165 983 9 996 DFRRQJI3VX1 $T=131040 69440 1 0 $X=130610 $Y=64320
X8754 1364 1362 165 1203 9 768 DFRRQJI3VX1 $T=131600 42560 0 0 $X=131170 $Y=41920
X8755 1364 1362 98 758 9 210 DFRRQJI3VX1 $T=148960 114240 0 180 $X=133410 $Y=109120
X8756 1364 1362 98 1198 15 234 DFRRQJI3VX1 $T=134960 141120 0 0 $X=134530 $Y=140480
X8757 1364 1362 98 221 15 229 DFRRQJI3VX1 $T=135520 159040 1 0 $X=135090 $Y=153920
X8758 1364 1362 98 5 15 266 DFRRQJI3VX1 $T=136080 141120 1 0 $X=135650 $Y=136000
X8759 1364 1362 178 1194 15 217 DFRRQJI3VX1 $T=136080 176960 0 0 $X=135650 $Y=176320
X8760 1364 1362 178 1195 15 993 DFRRQJI3VX1 $T=136640 194880 1 0 $X=136210 $Y=189760
X8761 1364 1362 233 6 15 1200 DFRRQJI3VX1 $T=138320 203840 0 0 $X=137890 $Y=203200
X8762 1364 1362 165 256 9 989 DFRRQJI3VX1 $T=160160 96320 1 180 $X=144610 $Y=95680
X8763 1364 1362 165 1305 9 1009 DFRRQJI3VX1 $T=145600 69440 0 0 $X=145170 $Y=68800
X8764 1364 1362 165 1006 9 997 DFRRQJI3VX1 $T=160720 105280 0 180 $X=145170 $Y=100160
X8765 1364 1362 165 238 9 1012 DFRRQJI3VX1 $T=147280 69440 1 0 $X=146850 $Y=64320
X8766 1364 1362 165 1205 9 251 DFRRQJI3VX1 $T=147840 42560 0 0 $X=147410 $Y=41920
X8767 1364 1362 165 1209 9 1000 DFRRQJI3VX1 $T=162960 51520 0 180 $X=147410 $Y=46400
X8768 1364 1362 165 1013 9 764 DFRRQJI3VX1 $T=162960 51520 1 180 $X=147410 $Y=50880
X8769 1364 1362 165 1208 9 763 DFRRQJI3VX1 $T=162960 60480 1 180 $X=147410 $Y=59840
X8770 1364 1362 98 773 15 249 DFRRQJI3VX1 $T=151200 159040 1 0 $X=150770 $Y=153920
X8771 1364 1362 98 1206 15 771 DFRRQJI3VX1 $T=166320 168000 1 180 $X=150770 $Y=167360
X8772 1364 1362 178 766 15 36 DFRRQJI3VX1 $T=166320 176960 1 180 $X=150770 $Y=176320
X8773 1364 1362 98 1207 15 236 DFRRQJI3VX1 $T=166880 150080 0 180 $X=151330 $Y=144960
X8774 1364 1362 233 265 15 1022 DFRRQJI3VX1 $T=151760 185920 1 0 $X=151330 $Y=180800
X8775 1364 1362 233 267 15 1017 DFRRQJI3VX1 $T=152320 185920 0 0 $X=151890 $Y=185280
X8776 1364 1362 233 268 15 295 DFRRQJI3VX1 $T=152320 194880 1 0 $X=151890 $Y=189760
X8777 1364 1362 233 1014 15 243 DFRRQJI3VX1 $T=170800 203840 1 180 $X=155250 $Y=203200
X8778 1364 1362 165 1018 9 776 DFRRQJI3VX1 $T=173600 105280 1 180 $X=158050 $Y=104640
X8779 1364 1362 165 1010 15 264 DFRRQJI3VX1 $T=159040 132160 0 0 $X=158610 $Y=131520
X8780 1364 1362 165 782 9 966 DFRRQJI3VX1 $T=175840 105280 0 180 $X=160290 $Y=100160
X8781 1364 1362 233 260 15 285 DFRRQJI3VX1 $T=160720 212800 0 0 $X=160290 $Y=212160
X8782 1364 1362 165 780 9 1016 DFRRQJI3VX1 $T=176960 96320 1 180 $X=161410 $Y=95680
X8783 1364 1362 165 255 9 1023 DFRRQJI3VX1 $T=163520 69440 1 0 $X=163090 $Y=64320
X8784 1364 1362 165 1210 9 252 DFRRQJI3VX1 $T=179200 42560 0 180 $X=163650 $Y=37440
X8785 1364 1362 165 1216 9 271 DFRRQJI3VX1 $T=179760 42560 1 180 $X=164210 $Y=41920
X8786 1364 1362 165 254 9 787 DFRRQJI3VX1 $T=164640 60480 1 0 $X=164210 $Y=55360
X8787 1364 1362 165 1212 9 263 DFRRQJI3VX1 $T=180320 51520 0 180 $X=164770 $Y=46400
X8788 1364 1362 165 792 9 1211 DFRRQJI3VX1 $T=165200 51520 0 0 $X=164770 $Y=50880
X8789 1364 1362 98 10 15 262 DFRRQJI3VX1 $T=181440 168000 0 180 $X=165890 $Y=162880
X8790 1364 1362 98 1021 15 279 DFRRQJI3VX1 $T=183120 159040 0 180 $X=167570 $Y=153920
X8791 1364 1362 165 1214 9 770 DFRRQJI3VX1 $T=188160 114240 0 180 $X=172610 $Y=109120
X8792 1364 1362 165 1028 15 278 DFRRQJI3VX1 $T=189840 132160 1 180 $X=174290 $Y=131520
X8793 1364 1362 165 1222 9 779 DFRRQJI3VX1 $T=190400 105280 1 180 $X=174850 $Y=104640
X8794 1364 1362 165 794 9 286 DFRRQJI3VX1 $T=190960 105280 0 180 $X=175410 $Y=100160
X8795 1364 1362 233 1027 15 311 DFRRQJI3VX1 $T=176960 212800 0 0 $X=176530 $Y=212160
X8796 1364 1362 165 1309 15 798 DFRRQJI3VX1 $T=193200 141120 1 180 $X=177650 $Y=140480
X8797 1364 1362 165 1220 9 296 DFRRQJI3VX1 $T=197120 42560 1 180 $X=181570 $Y=41920
X8798 1364 1362 165 1223 9 39 DFRRQJI3VX1 $T=197680 51520 0 180 $X=182130 $Y=46400
X8799 1364 1362 165 297 9 316 DFRRQJI3VX1 $T=182560 51520 0 0 $X=182130 $Y=50880
X8800 1364 1362 165 789 9 1036 DFRRQJI3VX1 $T=182560 60480 1 0 $X=182130 $Y=55360
X8801 1364 1362 165 336 9 277 DFRRQJI3VX1 $T=197680 123200 0 180 $X=182130 $Y=118080
X8802 1364 1362 320 1218 15 299 DFRRQJI3VX1 $T=197680 150080 0 180 $X=182130 $Y=144960
X8803 1364 1362 320 1224 15 292 DFRRQJI3VX1 $T=198240 150080 1 180 $X=182690 $Y=149440
X8804 1364 1362 165 1225 9 298 DFRRQJI3VX1 $T=198800 114240 1 180 $X=183250 $Y=113600
X8805 1364 1362 320 1333 15 340 DFRRQJI3VX1 $T=183680 159040 1 0 $X=183250 $Y=153920
X8806 1364 1362 320 1356 15 790 DFRRQJI3VX1 $T=184240 168000 1 0 $X=183810 $Y=162880
X8807 1364 1362 165 826 9 663 DFRRQJI3VX1 $T=203280 87360 1 180 $X=187730 $Y=86720
X8808 1364 1362 165 325 9 307 DFRRQJI3VX1 $T=203280 96320 0 180 $X=187730 $Y=91200
X8809 1364 1362 165 329 9 1030 DFRRQJI3VX1 $T=203280 114240 0 180 $X=187730 $Y=109120
X8810 1364 1362 165 1039 15 304 DFRRQJI3VX1 $T=203280 123200 1 180 $X=187730 $Y=122560
X8811 1364 1362 165 12 15 1217 DFRRQJI3VX1 $T=203280 132160 0 180 $X=187730 $Y=127040
X8812 1364 1362 339 1310 15 810 DFRRQJI3VX1 $T=192640 168000 0 0 $X=192210 $Y=167360
X8813 1364 1362 233 1228 15 328 DFRRQJI3VX1 $T=208320 212800 0 180 $X=192770 $Y=207680
X8814 1364 1362 320 321 15 1312 DFRRQJI3VX1 $T=198240 150080 1 0 $X=197810 $Y=144960
X8815 1364 1362 320 322 15 1157 DFRRQJI3VX1 $T=198240 150080 0 0 $X=197810 $Y=149440
X8816 1364 1362 320 1038 9 818 DFRRQJI3VX1 $T=199920 69440 1 0 $X=199490 $Y=64320
X8817 1364 1362 165 337 9 327 DFRRQJI3VX1 $T=215040 114240 1 180 $X=199490 $Y=113600
X8818 1364 1362 165 359 9 331 DFRRQJI3VX1 $T=215600 51520 0 180 $X=200050 $Y=46400
X8819 1364 1362 165 825 9 335 DFRRQJI3VX1 $T=215600 51520 1 180 $X=200050 $Y=50880
X8820 1364 1362 320 309 9 665 DFRRQJI3VX1 $T=201040 60480 0 0 $X=200610 $Y=59840
X8821 1364 1362 378 1311 9 346 DFRRQJI3VX1 $T=202720 60480 1 0 $X=202290 $Y=55360
X8822 1364 1362 822 1357 15 14 DFRRQJI3VX1 $T=204400 176960 0 0 $X=203970 $Y=176320
X8823 1364 1362 320 302 9 1043 DFRRQJI3VX1 $T=223440 69440 1 180 $X=207890 $Y=68800
X8824 1364 1362 233 1058 15 1045 DFRRQJI3VX1 $T=225680 212800 0 180 $X=210130 $Y=207680
X8825 1364 1362 320 811 15 814 DFRRQJI3VX1 $T=228480 141120 0 180 $X=212930 $Y=136000
X8826 1364 1362 320 1232 15 1048 DFRRQJI3VX1 $T=228480 141120 1 180 $X=212930 $Y=140480
X8827 1364 1362 320 1086 15 1020 DFRRQJI3VX1 $T=228480 150080 0 180 $X=212930 $Y=144960
X8828 1364 1362 819 392 15 1049 DFRRQJI3VX1 $T=228480 150080 1 180 $X=212930 $Y=149440
X8829 1364 1362 378 1314 15 1035 DFRRQJI3VX1 $T=228480 159040 1 180 $X=212930 $Y=158400
X8830 1364 1362 378 16 9 813 DFRRQJI3VX1 $T=226800 42560 1 0 $X=226370 $Y=37440
X8831 1364 1362 378 1237 9 381 DFRRQJI3VX1 $T=226800 51520 1 0 $X=226370 $Y=46400
X8832 1364 1362 378 1238 9 364 DFRRQJI3VX1 $T=226800 51520 0 0 $X=226370 $Y=50880
X8833 1364 1362 378 828 9 380 DFRRQJI3VX1 $T=226800 60480 1 0 $X=226370 $Y=55360
X8834 1364 1362 378 1056 9 1236 DFRRQJI3VX1 $T=226800 60480 0 0 $X=226370 $Y=59840
X8835 1364 1362 378 366 9 1064 DFRRQJI3VX1 $T=226800 69440 1 0 $X=226370 $Y=64320
X8836 1364 1362 379 1234 15 51 DFRRQJI3VX1 $T=226800 176960 0 0 $X=226370 $Y=176320
X8837 1364 1362 379 1315 15 839 DFRRQJI3VX1 $T=226800 185920 1 0 $X=226370 $Y=180800
X8838 1364 1362 379 1235 15 1065 DFRRQJI3VX1 $T=226800 194880 1 0 $X=226370 $Y=189760
X8839 1364 1362 379 827 15 1060 DFRRQJI3VX1 $T=226800 203840 0 0 $X=226370 $Y=203200
X8840 1364 1362 379 373 15 377 DFRRQJI3VX1 $T=229600 212800 1 0 $X=229170 $Y=207680
X8841 1364 1362 379 1062 15 837 DFRRQJI3VX1 $T=230720 159040 1 0 $X=230290 $Y=153920
X8842 1364 1362 379 667 15 383 DFRRQJI3VX1 $T=231280 150080 0 0 $X=230850 $Y=149440
X8843 1364 1362 379 387 15 1073 DFRRQJI3VX1 $T=232960 141120 0 0 $X=232530 $Y=140480
X8844 1364 1362 395 375 9 396 DFRRQJI3VX1 $T=236320 114240 1 0 $X=235890 $Y=109120
X8845 1364 1362 391 823 15 668 DFRRQJI3VX1 $T=236880 132160 0 0 $X=236450 $Y=131520
X8846 1364 1362 378 1242 9 399 DFRRQJI3VX1 $T=239120 42560 0 0 $X=238690 $Y=41920
X8847 1364 1362 395 382 15 1247 DFRRQJI3VX1 $T=240240 123200 0 0 $X=239810 $Y=122560
X8848 1364 1362 395 1074 15 846 DFRRQJI3VX1 $T=240240 132160 1 0 $X=239810 $Y=127040
X8849 1364 1362 379 1318 15 843 DFRRQJI3VX1 $T=240240 203840 1 0 $X=239810 $Y=198720
X8850 1364 1362 378 1245 9 409 DFRRQJI3VX1 $T=241920 42560 1 0 $X=241490 $Y=37440
X8851 1364 1362 378 1249 9 1066 DFRRQJI3VX1 $T=257040 51520 0 180 $X=241490 $Y=46400
X8852 1364 1362 378 829 9 1077 DFRRQJI3VX1 $T=241920 51520 0 0 $X=241490 $Y=50880
X8853 1364 1362 378 1079 9 832 DFRRQJI3VX1 $T=257040 60480 0 180 $X=241490 $Y=55360
X8854 1364 1362 378 371 9 1067 DFRRQJI3VX1 $T=257040 60480 1 180 $X=241490 $Y=59840
X8855 1364 1362 378 830 9 835 DFRRQJI3VX1 $T=257040 69440 0 180 $X=241490 $Y=64320
X8856 1364 1362 379 1319 15 393 DFRRQJI3VX1 $T=259840 203840 1 180 $X=244290 $Y=203200
X8857 1364 1362 379 1257 15 397 DFRRQJI3VX1 $T=261520 150080 1 180 $X=245970 $Y=149440
X8858 1364 1362 379 1081 15 390 DFRRQJI3VX1 $T=261520 159040 0 180 $X=245970 $Y=153920
X8859 1364 1362 379 1248 15 417 DFRRQJI3VX1 $T=249200 212800 1 0 $X=248770 $Y=207680
X8860 1364 1362 379 403 15 1243 DFRRQJI3VX1 $T=265440 150080 0 180 $X=249890 $Y=144960
X8861 1364 1362 378 1078 9 1254 DFRRQJI3VX1 $T=252000 69440 0 0 $X=251570 $Y=68800
X8862 1364 1362 395 1091 15 414 DFRRQJI3VX1 $T=272160 132160 0 180 $X=256610 $Y=127040
X8863 1364 1362 378 1258 9 413 DFRRQJI3VX1 $T=272720 51520 0 180 $X=257170 $Y=46400
X8864 1364 1362 378 1261 9 437 DFRRQJI3VX1 $T=257600 51520 0 0 $X=257170 $Y=50880
X8865 1364 1362 378 450 9 442 DFRRQJI3VX1 $T=257600 60480 0 0 $X=257170 $Y=59840
X8866 1364 1362 378 847 9 669 DFRRQJI3VX1 $T=272720 69440 0 180 $X=257170 $Y=64320
X8867 1364 1362 378 1253 9 441 DFRRQJI3VX1 $T=258160 60480 1 0 $X=257730 $Y=55360
X8868 1364 1362 395 451 15 1259 DFRRQJI3VX1 $T=259280 123200 0 0 $X=258850 $Y=122560
X8869 1364 1362 395 386 9 1088 DFRRQJI3VX1 $T=259840 123200 1 0 $X=259410 $Y=118080
X8870 1364 1362 379 1090 15 432 DFRRQJI3VX1 $T=276080 159040 1 180 $X=260530 $Y=158400
X8871 1364 1362 379 1256 15 428 DFRRQJI3VX1 $T=276080 203840 1 180 $X=260530 $Y=203200
X8872 1364 1362 379 1262 15 1251 DFRRQJI3VX1 $T=277200 159040 0 180 $X=261650 $Y=153920
X8873 1364 1362 379 443 15 420 DFRRQJI3VX1 $T=277760 150080 1 180 $X=262210 $Y=149440
X8874 1364 1362 378 427 9 430 DFRRQJI3VX1 $T=282240 69440 1 180 $X=266690 $Y=68800
X8875 1364 1362 378 1094 9 453 DFRRQJI3VX1 $T=291200 51520 0 180 $X=275650 $Y=46400
X8876 1364 1362 378 1266 9 458 DFRRQJI3VX1 $T=291200 51520 1 180 $X=275650 $Y=50880
X8877 1364 1362 378 1097 9 457 DFRRQJI3VX1 $T=291200 60480 0 180 $X=275650 $Y=55360
X8878 1364 1362 378 444 9 1095 DFRRQJI3VX1 $T=276080 60480 0 0 $X=275650 $Y=59840
X8879 1364 1362 378 1260 9 867 DFRRQJI3VX1 $T=276080 69440 1 0 $X=275650 $Y=64320
X8880 1364 1362 378 454 9 670 DFRRQJI3VX1 $T=276640 96320 1 0 $X=276210 $Y=91200
X8881 1364 1362 395 18 15 45 DFRRQJI3VX1 $T=291760 123200 0 180 $X=276210 $Y=118080
X8882 1364 1362 395 863 15 473 DFRRQJI3VX1 $T=277200 123200 0 0 $X=276770 $Y=122560
X8883 1364 1362 379 860 15 17 DFRRQJI3VX1 $T=292320 194880 1 180 $X=276770 $Y=194240
X8884 1364 1362 395 481 15 870 DFRRQJI3VX1 $T=277760 159040 0 0 $X=277330 $Y=158400
X8885 1364 1362 395 461 15 476 DFRRQJI3VX1 $T=278320 159040 1 0 $X=277890 $Y=153920
X8886 1364 1362 379 1267 15 459 DFRRQJI3VX1 $T=293440 168000 0 180 $X=277890 $Y=162880
X8887 1364 1362 379 868 15 861 DFRRQJI3VX1 $T=295120 176960 0 180 $X=279570 $Y=171840
X8888 1364 1362 379 864 15 447 DFRRQJI3VX1 $T=295120 194880 0 180 $X=279570 $Y=189760
X8889 1364 1362 395 508 19 490 DFRRQJI3VX1 $T=292320 150080 0 0 $X=291890 $Y=149440
X8890 1364 1362 378 1269 9 475 DFRRQJI3VX1 $T=309120 51520 0 180 $X=293570 $Y=46400
X8891 1364 1362 378 1274 9 872 DFRRQJI3VX1 $T=309120 51520 1 180 $X=293570 $Y=50880
X8892 1364 1362 378 1271 9 474 DFRRQJI3VX1 $T=309120 60480 0 180 $X=293570 $Y=55360
X8893 1364 1362 378 1100 9 1268 DFRRQJI3VX1 $T=294000 60480 0 0 $X=293570 $Y=59840
X8894 1364 1362 378 501 9 671 DFRRQJI3VX1 $T=294000 69440 1 0 $X=293570 $Y=64320
X8895 1364 1362 395 495 19 361 DFRRQJI3VX1 $T=309120 159040 1 180 $X=293570 $Y=158400
X8896 1364 1362 378 505 9 672 DFRRQJI3VX1 $T=294560 78400 1 0 $X=294130 $Y=73280
X8897 1364 1362 378 1272 9 1098 DFRRQJI3VX1 $T=310240 42560 0 180 $X=294690 $Y=37440
X8898 1364 1362 378 506 9 494 DFRRQJI3VX1 $T=295120 69440 0 0 $X=294690 $Y=68800
X8899 1364 1362 533 875 33 498 DFRRQJI3VX1 $T=297360 212800 1 0 $X=296930 $Y=207680
X8900 1364 1362 395 873 19 521 DFRRQJI3VX1 $T=307440 150080 0 0 $X=307010 $Y=149440
X8901 1364 1362 378 1278 19 503 DFRRQJI3VX1 $T=326480 51520 0 180 $X=310930 $Y=46400
X8902 1364 1362 378 1276 19 55 DFRRQJI3VX1 $T=326480 51520 1 180 $X=310930 $Y=50880
X8903 1364 1362 378 540 19 513 DFRRQJI3VX1 $T=326480 60480 0 180 $X=310930 $Y=55360
X8904 1364 1362 378 551 19 1103 DFRRQJI3VX1 $T=326480 69440 0 180 $X=310930 $Y=64320
X8905 1364 1362 395 1322 19 534 DFRRQJI3VX1 $T=311360 185920 1 0 $X=310930 $Y=180800
X8906 1364 1362 378 539 19 1109 DFRRQJI3VX1 $T=311920 42560 1 0 $X=311490 $Y=37440
X8907 1364 1362 378 550 19 674 DFRRQJI3VX1 $T=327040 60480 1 180 $X=311490 $Y=59840
X8908 1364 1362 378 546 19 1280 DFRRQJI3VX1 $T=311920 69440 0 0 $X=311490 $Y=68800
X8909 1364 1362 378 514 19 673 DFRRQJI3VX1 $T=311920 78400 1 0 $X=311490 $Y=73280
X8910 1364 1362 395 1102 19 532 DFRRQJI3VX1 $T=311920 185920 0 0 $X=311490 $Y=185280
X8911 1364 1362 533 1106 33 502 DFRRQJI3VX1 $T=327600 203840 1 180 $X=312050 $Y=203200
X8912 1364 1362 533 512 33 519 DFRRQJI3VX1 $T=314720 203840 1 0 $X=314290 $Y=198720
X8913 1364 1362 395 1279 19 893 DFRRQJI3VX1 $T=322000 132160 1 0 $X=321570 $Y=127040
X8914 1364 1362 395 515 19 894 DFRRQJI3VX1 $T=322000 132160 0 0 $X=321570 $Y=131520
X8915 1364 1362 395 883 19 1285 DFRRQJI3VX1 $T=322000 141120 1 0 $X=321570 $Y=136000
X8916 1364 1362 395 1324 19 528 DFRRQJI3VX1 $T=337120 150080 0 180 $X=321570 $Y=144960
X8917 1364 1362 395 1323 19 553 DFRRQJI3VX1 $T=322000 159040 1 0 $X=321570 $Y=153920
X8918 1364 1362 395 516 19 679 DFRRQJI3VX1 $T=322560 141120 0 0 $X=322130 $Y=140480
X8919 1364 1362 395 517 19 895 DFRRQJI3VX1 $T=322560 150080 0 0 $X=322130 $Y=149440
X8920 1364 1362 395 1275 19 523 DFRRQJI3VX1 $T=338240 159040 1 180 $X=322690 $Y=158400
X8921 1364 1362 378 1288 19 535 DFRRQJI3VX1 $T=342720 51520 0 180 $X=327170 $Y=46400
X8922 1364 1362 378 569 19 537 DFRRQJI3VX1 $T=342720 51520 1 180 $X=327170 $Y=50880
X8923 1364 1362 378 574 19 1114 DFRRQJI3VX1 $T=328160 60480 1 0 $X=327730 $Y=55360
X8924 1364 1362 378 573 19 675 DFRRQJI3VX1 $T=328160 69440 1 0 $X=327730 $Y=64320
X8925 1364 1362 395 548 19 544 DFRRQJI3VX1 $T=329280 185920 0 0 $X=328850 $Y=185280
X8926 1364 1362 395 1284 19 57 DFRRQJI3VX1 $T=329840 194880 0 0 $X=329410 $Y=194240
X8927 1364 1362 533 1345 33 676 DFRRQJI3VX1 $T=336000 203840 0 0 $X=335570 $Y=203200
X8928 1364 1362 395 20 19 939 DFRRQJI3VX1 $T=355040 132160 0 180 $X=339490 $Y=127040
X8929 1364 1362 395 1289 19 552 DFRRQJI3VX1 $T=355040 150080 1 180 $X=339490 $Y=149440
X8930 1364 1362 395 564 19 561 DFRRQJI3VX1 $T=355040 159040 0 180 $X=339490 $Y=153920
X8931 1364 1362 395 541 19 677 DFRRQJI3VX1 $T=355600 132160 1 180 $X=340050 $Y=131520
X8932 1364 1362 395 1132 19 619 DFRRQJI3VX1 $T=355600 141120 0 180 $X=340050 $Y=136000
X8933 1364 1362 395 1125 19 554 DFRRQJI3VX1 $T=355600 150080 0 180 $X=340050 $Y=144960
X8934 1364 1362 395 1283 19 560 DFRRQJI3VX1 $T=356720 42560 1 180 $X=341170 $Y=41920
X8935 1364 1362 395 580 19 1113 DFRRQJI3VX1 $T=356720 60480 1 180 $X=341170 $Y=59840
X8936 1364 1362 395 1118 19 1128 DFRRQJI3VX1 $T=355040 51520 0 0 $X=354610 $Y=50880
X8937 1364 1362 22 907 19 589 DFRRQJI3VX1 $T=355040 69440 1 0 $X=354610 $Y=64320
X8938 1364 1362 22 576 19 581 DFRRQJI3VX1 $T=355040 194880 1 0 $X=354610 $Y=189760
X8939 1364 1362 22 1290 19 575 DFRRQJI3VX1 $T=355040 194880 0 0 $X=354610 $Y=194240
X8940 1364 1362 22 601 19 915 DFRRQJI3VX1 $T=357280 150080 0 0 $X=356850 $Y=149440
X8941 1364 1362 22 602 19 940 DFRRQJI3VX1 $T=357840 159040 1 0 $X=357410 $Y=153920
X8942 1364 1362 22 1293 19 1295 DFRRQJI3VX1 $T=358400 141120 1 0 $X=357970 $Y=136000
X8943 1364 1362 22 1130 19 607 DFRRQJI3VX1 $T=358400 141120 0 0 $X=357970 $Y=140480
X8944 1364 1362 22 596 19 905 DFRRQJI3VX1 $T=358400 159040 0 0 $X=357970 $Y=158400
X8945 1364 1362 22 1129 19 1119 DFRRQJI3VX1 $T=358400 168000 1 0 $X=357970 $Y=162880
X8946 1364 1362 22 599 19 604 DFRRQJI3VX1 $T=358960 132160 0 0 $X=358530 $Y=131520
X8947 1364 1362 395 1296 19 678 DFRRQJI3VX1 $T=377440 42560 1 180 $X=361890 $Y=41920
X8948 1364 1362 22 1136 19 1133 DFRRQJI3VX1 $T=362320 60480 0 0 $X=361890 $Y=59840
X8949 1364 1362 395 916 19 61 DFRRQJI3VX1 $T=378000 51520 0 180 $X=362450 $Y=46400
X8950 1364 1362 22 600 19 1134 DFRRQJI3VX1 $T=362880 60480 1 0 $X=362450 $Y=55360
X8951 1364 1362 22 605 19 587 DFRRQJI3VX1 $T=380800 176960 1 180 $X=365250 $Y=176320
X8952 1364 1362 22 1137 19 680 DFRRQJI3VX1 $T=381360 176960 0 180 $X=365810 $Y=171840
X8953 1364 1362 22 918 19 591 DFRRQJI3VX1 $T=388640 150080 1 180 $X=373090 $Y=149440
X8954 1364 1362 22 62 19 595 DFRRQJI3VX1 $T=394800 51520 0 180 $X=379250 $Y=46400
X8955 1364 1362 22 1328 19 592 DFRRQJI3VX1 $T=395360 42560 0 180 $X=379810 $Y=37440
X8956 1364 1362 22 1298 19 598 DFRRQJI3VX1 $T=395360 42560 1 180 $X=379810 $Y=41920
X8957 1364 1362 22 1145 19 590 DFRRQJI3VX1 $T=395360 51520 1 180 $X=379810 $Y=50880
X8958 1364 1362 22 682 19 922 DFRRQJI3VX1 $T=380240 60480 1 0 $X=379810 $Y=55360
X8959 1364 1362 22 681 19 632 DFRRQJI3VX1 $T=380240 60480 0 0 $X=379810 $Y=59840
X8960 1364 1362 22 917 19 923 DFRRQJI3VX1 $T=380240 69440 1 0 $X=379810 $Y=64320
X8961 1364 1362 22 611 19 1144 DFRRQJI3VX1 $T=380240 69440 0 0 $X=379810 $Y=68800
X8962 1364 1362 22 929 19 628 DFRRQJI3VX1 $T=408800 150080 1 180 $X=393250 $Y=149440
X8963 1364 1362 22 924 19 626 DFRRQJI3VX1 $T=409920 132160 0 180 $X=394370 $Y=127040
X8964 1364 1362 22 645 19 640 DFRRQJI3VX1 $T=413280 42560 0 180 $X=397730 $Y=37440
X8965 1364 1362 22 646 19 930 DFRRQJI3VX1 $T=413280 42560 1 180 $X=397730 $Y=41920
X8966 1364 1362 22 647 19 637 DFRRQJI3VX1 $T=413280 51520 0 180 $X=397730 $Y=46400
X8967 1364 1362 22 648 19 635 DFRRQJI3VX1 $T=413280 51520 1 180 $X=397730 $Y=50880
X8968 1364 1362 22 638 19 684 DFRRQJI3VX1 $T=398160 60480 1 0 $X=397730 $Y=55360
X8969 1364 1362 22 1150 19 683 DFRRQJI3VX1 $T=398160 60480 0 0 $X=397730 $Y=59840
X8970 1364 1362 22 23 19 934 DFRRQJI3VX1 $T=398160 69440 1 0 $X=397730 $Y=64320
X8971 1364 1362 22 24 19 644 DFRRQJI3VX1 $T=398160 69440 0 0 $X=397730 $Y=68800
X8972 1364 1362 22 25 19 462 DFRRQJI3VX1 $T=398160 105280 1 0 $X=397730 $Y=100160
X8973 1364 1362 71 85 INJI3VX1 $T=42000 159040 1 0 $X=41570 $Y=153920
X8974 1364 1362 80 948 INJI3VX1 $T=42560 176960 0 0 $X=42130 $Y=176320
X8975 1364 1362 91 951 INJI3VX1 $T=50960 176960 0 0 $X=50530 $Y=176320
X8976 1364 1362 654 111 INJI3VX1 $T=63840 194880 1 0 $X=63410 $Y=189760
X8977 1364 1362 152 1026 INJI3VX1 $T=181440 150080 0 0 $X=181010 $Y=149440
X8978 1364 1362 45 140 INJI3VX1 $T=202720 176960 0 0 $X=202290 $Y=176320
X8979 1364 1362 152 1061 INJI3VX1 $T=231840 176960 1 0 $X=231410 $Y=171840
X8980 1364 1362 1061 379 INJI3VX1 $T=233520 168000 0 0 $X=233090 $Y=167360
X8981 1364 1362 377 1063 INJI3VX1 $T=238560 203840 1 0 $X=238130 $Y=198720
X8982 1364 1362 843 844 INJI3VX1 $T=247520 185920 0 0 $X=247090 $Y=185280
X8983 1364 1362 41 533 INJI3VX1 $T=309120 203840 0 0 $X=308690 $Y=203200
X8984 1364 1362 626 613 INJI3VX1 $T=392560 132160 1 0 $X=392130 $Y=127040
X8985 1364 1362 1026 98 INJI3VX2 $T=180320 150080 1 0 $X=179890 $Y=144960
X8986 1364 1362 125 DAC<1> BUJI3VX12 $T=69440 24640 0 180 $X=56690 $Y=19520
X8987 1364 1362 725 DAC<2> BUJI3VX12 $T=77840 24640 1 180 $X=65090 $Y=24000
X8988 1364 1362 726 DAC<3> BUJI3VX12 $T=82880 24640 0 180 $X=70130 $Y=19520
X8989 1364 1362 78 81 65 943 69 ON22JI3VX1 $T=33600 159040 0 180 $X=28690 $Y=153920
X8990 1364 1362 75 945 1395 74 68 ON22JI3VX1 $T=36400 168000 1 180 $X=31490 $Y=167360
X8991 1364 1362 691 79 696 948 693 ON22JI3VX1 $T=40320 168000 1 0 $X=39890 $Y=162880
X8992 1364 1362 653 1390 1168 96 1167 ON22JI3VX1 $T=58800 185920 1 180 $X=53890 $Y=185280
X8993 1364 1362 706 111 1172 1171 1394 ON22JI3VX1 $T=63280 168000 0 0 $X=62850 $Y=167360
X8994 1364 1362 1171 139 119 96 124 ON22JI3VX1 $T=71680 194880 0 180 $X=66770 $Y=189760
X8995 1364 1362 1317 423 1315 1070 385 ON22JI3VX1 $T=246400 185920 0 180 $X=241490 $Y=180800
X8996 1364 1362 400 423 1319 1246 410 ON22JI3VX1 $T=251440 194880 1 0 $X=251010 $Y=189760
X8997 1364 1362 432 431 849 1083 1251 ON22JI3VX1 $T=267680 185920 1 180 $X=262770 $Y=185280
X8998 1364 1362 528 884 507 1107 523 ON22JI3VX1 $T=319760 159040 1 180 $X=314850 $Y=158400
X8999 1364 1362 544 556 1286 900 57 ON22JI3VX1 $T=344960 185920 0 180 $X=340050 $Y=180800
X9000 1364 1362 587 1123 547 21 1119 ON22JI3VX1 $T=364560 168000 1 180 $X=359650 $Y=167360
X9001 1364 1362 636 633 621 617 639 ON22JI3VX1 $T=392560 114240 0 180 $X=387650 $Y=109120
X9002 1364 1362 641 925 929 941 628 ON22JI3VX1 $T=398720 159040 1 0 $X=398290 $Y=153920
X9003 1364 1362 1219 324 802 42 333 AN31JI3VX1 $T=195440 185920 0 0 $X=195010 $Y=185280
X9004 1364 1362 425 1084 845 1255 446 AN31JI3VX1 $T=264320 168000 0 0 $X=263890 $Y=167360
X9005 1364 1362 1396 1273 1343 492 1270 AN31JI3VX1 $T=313040 168000 0 180 $X=308690 $Y=162880
X9006 1364 1362 1353 121 1397 1172 NO3JI3VX0 $T=63840 176960 1 0 $X=63410 $Y=171840
X9007 1364 1362 1380 1376 1068 389 NO3JI3VX0 $T=246400 159040 0 0 $X=245970 $Y=158400
X9008 1364 1362 477 485 1398 493 NO3JI3VX0 $T=295120 212800 0 0 $X=294690 $Y=212160
X9009 1364 1362 140 530 54 877 NO3JI3VX0 $T=305200 176960 0 0 $X=304770 $Y=176320
X9010 1364 1362 313 319 115 809 343 OR4JI3VX2 $T=194320 24640 0 0 $X=193890 $Y=24000
X9011 1364 1362 1152 215 35 208 HAJI3VX1 $T=138320 203840 1 180 $X=130050 $Y=203200
X9012 1364 1362 1399 215 243 767 HAJI3VX1 $T=158480 212800 0 180 $X=150210 $Y=207680
X9013 1364 1362 785 272 1022 276 HAJI3VX1 $T=175840 185920 0 180 $X=167570 $Y=180800
X9014 1364 1362 282 1019 285 786 HAJI3VX1 $T=173600 203840 0 0 $X=173170 $Y=203200
X9015 1364 1362 1400 1017 276 293 HAJI3VX1 $T=175280 185920 0 0 $X=174850 $Y=185280
X9016 1364 1362 796 311 786 46 HAJI3VX1 $T=186480 203840 0 0 $X=186050 $Y=203200
X9017 1364 1362 418 417 1401 412 HAJI3VX1 $T=262080 194880 1 180 $X=253810 $Y=194240
X9018 1364 1362 424 428 412 421 HAJI3VX1 $T=267680 203840 0 180 $X=259410 $Y=198720
X9019 1364 1362 512 519 885 509 HAJI3VX1 $T=316960 212800 1 0 $X=316530 $Y=207680
X9020 1364 1362 526 1096 532 1281 HAJI3VX1 $T=322000 176960 0 0 $X=321570 $Y=176320
X9021 1364 1362 1111 536 1402 885 HAJI3VX1 $T=329840 212800 0 0 $X=329410 $Y=212160
X9022 1364 1362 1120 575 899 1122 HAJI3VX1 $T=351680 176960 1 180 $X=343410 $Y=176320
X9023 1364 1362 1252 374 DLY4JI3VX1 $T=252000 212800 0 0 $X=251570 $Y=212160
X9024 1364 1362 702 1374 94 NO2I1JI3VX1 $T=50400 150080 0 0 $X=49970 $Y=149440
X9025 1364 1362 770 230 229 NO2I1JI3VX1 $T=143360 123200 0 0 $X=142930 $Y=122560
X9026 1364 1362 779 247 249 NO2I1JI3VX1 $T=166320 132160 0 180 $X=162530 $Y=127040
X9027 1364 1362 299 40 1017 NO2I1JI3VX1 $T=184240 185920 0 0 $X=183810 $Y=185280
X9028 1364 1362 1017 1034 299 NO2I1JI3VX1 $T=187600 185920 0 0 $X=187170 $Y=185280
X9029 1364 1362 308 11 310 NO2I1JI3VX1 $T=187600 203840 1 0 $X=187170 $Y=198720
X9030 1364 1362 340 323 361 NO2I1JI3VX1 $T=197680 176960 1 0 $X=197250 $Y=171840
X9031 1364 1362 808 231 47 NO2I1JI3VX1 $T=202720 168000 0 180 $X=198930 $Y=162880
X9032 1364 1362 806 353 347 NO2I1JI3VX1 $T=210000 159040 0 180 $X=206210 $Y=153920
X9033 1364 1362 1060 13 361 NO2I1JI3VX1 $T=219520 194880 1 180 $X=215730 $Y=194240
X9034 1364 1362 361 1057 1060 NO2I1JI3VX1 $T=235200 194880 1 180 $X=231410 $Y=194240
X9035 1364 1362 840 402 404 NO2I1JI3VX1 $T=249760 168000 1 0 $X=249330 $Y=162880
X9036 1364 1362 861 446 447 NO2I1JI3VX1 $T=278320 176960 0 180 $X=274530 $Y=171840
X9037 1364 1362 456 857 459 NO2I1JI3VX1 $T=280560 168000 1 180 $X=276770 $Y=167360
X9038 1364 1362 485 1104 496 NO2I1JI3VX1 $T=306880 123200 0 0 $X=306450 $Y=122560
X9039 1364 1362 525 1344 523 NO2I1JI3VX1 $T=332640 168000 0 180 $X=328850 $Y=162880
X9040 1364 1362 552 543 544 NO2I1JI3VX1 $T=337120 176960 0 180 $X=333330 $Y=171840
X9041 1364 1362 544 881 552 NO2I1JI3VX1 $T=338800 168000 1 180 $X=335010 $Y=167360
X9042 1364 1362 70 1395 87 68 685 AO22JI3VX1 $T=31360 168000 1 180 $X=25890 $Y=167360
X9043 1364 1362 88 70 80 140 67 AO22JI3VX1 $T=44240 185920 1 180 $X=38770 $Y=185280
X9044 1364 1362 701 70 953 140 89 AO22JI3VX1 $T=50960 185920 1 180 $X=45490 $Y=185280
X9045 1364 1362 721 245 148 143 141 AO22JI3VX1 $T=86800 42560 0 180 $X=81330 $Y=37440
X9046 1364 1362 157 245 148 727 142 AO22JI3VX1 $T=89040 33600 0 180 $X=83570 $Y=28480
X9047 1364 1362 724 245 148 709 365 AO22JI3VX1 $T=95200 33600 0 180 $X=89730 $Y=28480
X9048 1364 1362 153 245 148 733 388 AO22JI3VX1 $T=103040 33600 0 0 $X=102610 $Y=32960
X9049 1364 1362 164 245 148 163 422 AO22JI3VX1 $T=109760 33600 0 0 $X=109330 $Y=32960
X9050 1364 1362 174 245 148 167 338 AO22JI3VX1 $T=112000 33600 1 0 $X=111570 $Y=28480
X9051 1364 1362 987 240 237 749 195 AO22JI3VX1 $T=130480 203840 1 180 $X=125010 $Y=203200
X9052 1364 1362 192 245 148 752 342 AO22JI3VX1 $T=126560 24640 0 0 $X=126130 $Y=24000
X9053 1364 1362 754 240 237 223 189 AO22JI3VX1 $T=131600 141120 1 180 $X=126130 $Y=140480
X9054 1364 1362 755 240 237 979 190 AO22JI3VX1 $T=132160 159040 0 180 $X=126690 $Y=153920
X9055 1364 1362 976 240 237 980 194 AO22JI3VX1 $T=132160 185920 0 180 $X=126690 $Y=180800
X9056 1364 1362 991 240 237 978 660 AO22JI3VX1 $T=133840 194880 1 180 $X=128370 $Y=194240
X9057 1364 1362 197 240 237 981 1191 AO22JI3VX1 $T=129360 168000 1 0 $X=128930 $Y=162880
X9058 1364 1362 1152 240 237 35 1197 AO22JI3VX1 $T=137760 212800 1 0 $X=137330 $Y=207680
X9059 1364 1362 765 246 43 217 1194 AO22JI3VX1 $T=146160 168000 1 180 $X=140690 $Y=167360
X9060 1364 1362 219 246 43 36 766 AO22JI3VX1 $T=141680 185920 1 0 $X=141250 $Y=180800
X9061 1364 1362 1004 246 43 993 1195 AO22JI3VX1 $T=146720 194880 1 180 $X=141250 $Y=194240
X9062 1364 1362 205 245 148 214 348 AO22JI3VX1 $T=142240 33600 0 0 $X=141810 $Y=32960
X9063 1364 1362 992 246 43 1200 6 AO22JI3VX1 $T=143360 212800 1 0 $X=142930 $Y=207680
X9064 1364 1362 1202 246 43 229 221 AO22JI3VX1 $T=150640 159040 1 180 $X=145170 $Y=158400
X9065 1364 1362 226 245 148 768 357 AO22JI3VX1 $T=148960 24640 0 0 $X=148530 $Y=24000
X9066 1364 1362 235 246 43 249 773 AO22JI3VX1 $T=150640 159040 0 0 $X=150210 $Y=158400
X9067 1364 1362 240 778 237 236 1207 AO22JI3VX1 $T=155120 141120 1 0 $X=154690 $Y=136000
X9068 1364 1362 763 245 148 1000 330 AO22JI3VX1 $T=156240 33600 0 0 $X=155810 $Y=32960
X9069 1364 1362 246 259 43 771 1206 AO22JI3VX1 $T=163520 159040 1 180 $X=158050 $Y=158400
X9070 1364 1362 240 1306 237 264 1010 AO22JI3VX1 $T=165760 141120 0 180 $X=160290 $Y=136000
X9071 1364 1362 1399 246 43 269 1014 AO22JI3VX1 $T=160720 212800 1 0 $X=160290 $Y=207680
X9072 1364 1362 252 245 148 251 398 AO22JI3VX1 $T=163520 33600 1 0 $X=163090 $Y=28480
X9073 1364 1362 246 781 43 262 10 AO22JI3VX1 $T=166880 159040 0 0 $X=166450 $Y=158400
X9074 1364 1362 785 240 237 1022 265 AO22JI3VX1 $T=174160 176960 1 180 $X=168690 $Y=176320
X9075 1364 1362 1400 240 237 1017 267 AO22JI3VX1 $T=174160 185920 1 180 $X=168690 $Y=185280
X9076 1364 1362 1403 240 237 295 268 AO22JI3VX1 $T=174160 194880 0 180 $X=168690 $Y=189760
X9077 1364 1362 282 246 43 285 260 AO22JI3VX1 $T=174160 212800 0 180 $X=168690 $Y=207680
X9078 1364 1362 271 245 148 263 283 AO22JI3VX1 $T=170240 24640 0 0 $X=169810 $Y=24000
X9079 1364 1362 246 1331 43 279 1021 AO22JI3VX1 $T=181440 159040 1 180 $X=175970 $Y=158400
X9080 1364 1362 240 788 237 278 1028 AO22JI3VX1 $T=180320 141120 1 0 $X=179890 $Y=136000
X9081 1364 1362 796 246 43 311 1027 AO22JI3VX1 $T=187040 212800 0 180 $X=181570 $Y=207680
X9082 1364 1362 296 245 148 39 439 AO22JI3VX1 $T=187040 33600 0 0 $X=186610 $Y=32960
X9083 1364 1362 1404 246 43 328 1228 AO22JI3VX1 $T=201040 203840 0 0 $X=200610 $Y=203200
X9084 1364 1362 335 245 148 331 354 AO22JI3VX1 $T=205520 42560 1 0 $X=205090 $Y=37440
X9085 1364 1362 418 1153 1239 417 1248 AO22JI3VX1 $T=260960 194880 0 180 $X=255490 $Y=189760
X9086 1364 1362 416 411 849 854 1085 AO22JI3VX1 $T=259840 176960 0 0 $X=259410 $Y=176320
X9087 1364 1362 424 1153 1239 428 1256 AO22JI3VX1 $T=262640 194880 0 0 $X=262210 $Y=194240
X9088 1364 1362 413 426 384 437 579 AO22JI3VX1 $T=266560 33600 1 0 $X=266130 $Y=28480
X9089 1364 1362 448 1153 1239 17 860 AO22JI3VX1 $T=270480 194880 0 0 $X=270050 $Y=194240
X9090 1364 1362 474 426 384 475 876 AO22JI3VX1 $T=299040 33600 1 0 $X=298610 $Y=28480
X9091 1364 1362 526 530 877 532 1102 AO22JI3VX1 $T=314720 194880 0 180 $X=309250 $Y=189760
X9092 1364 1362 522 530 877 534 1322 AO22JI3VX1 $T=320880 176960 1 180 $X=315410 $Y=176320
X9093 1364 1362 513 426 384 55 577 AO22JI3VX1 $T=320320 33600 0 0 $X=319890 $Y=32960
X9094 1364 1362 503 426 384 1109 887 AO22JI3VX1 $T=320880 33600 1 0 $X=320450 $Y=28480
X9095 1364 1362 57 542 530 1286 1284 AO22JI3VX1 $T=341600 194880 0 180 $X=336130 $Y=189760
X9096 1364 1362 1120 530 877 575 1290 AO22JI3VX1 $T=352240 185920 1 180 $X=346770 $Y=185280
X9097 1364 1362 115 pulse_active BUJI3VX6 $T=55440 24640 0 0 $X=55010 $Y=24000
X9098 1364 1362 723 33 BUJI3VX6 $T=77280 123200 0 0 $X=76850 $Y=122560
X9099 1364 1362 1405 395 BUJI3VX6 $T=285600 132160 0 0 $X=285170 $Y=131520
X9100 1364 1362 591 384 BUJI3VX6 $T=373520 150080 1 0 $X=373090 $Y=144960
X9101 1364 1362 71 69 81 942 1406 ON31JI3VX1 $T=32480 150080 1 180 $X=27570 $Y=149440
X9102 1364 1362 75 946 96 66 1407 ON31JI3VX1 $T=36960 176960 1 180 $X=32050 $Y=176320
X9103 1364 1362 654 118 96 3 710 ON31JI3VX1 $T=63840 194880 0 180 $X=58930 $Y=189760
X9104 1364 1362 790 290 288 1356 1332 ON31JI3VX1 $T=180320 168000 0 0 $X=179890 $Y=167360
X9105 1364 1362 1045 349 1335 1058 1231 ON31JI3VX1 $T=211120 203840 0 0 $X=210690 $Y=203200
X9106 1364 1362 843 1241 423 1318 1240 ON31JI3VX1 $T=249760 194880 1 180 $X=244850 $Y=194240
X9107 1364 1362 447 855 423 864 862 ON31JI3VX1 $T=274400 194880 1 0 $X=273970 $Y=189760
X9108 1364 1362 1281 1277 1344 524 529 ON31JI3VX1 $T=328720 168000 1 180 $X=323810 $Y=167360
X9109 1364 1362 544 545 903 548 891 ON31JI3VX1 $T=331520 185920 1 0 $X=331090 $Y=180800
X9110 1364 1362 581 902 903 576 586 ON31JI3VX1 $T=347200 194880 1 0 $X=346770 $Y=189760
X9111 1364 1362 626 1297 63 924 1408 ON31JI3VX1 $T=392000 123200 1 0 $X=391570 $Y=118080
X9112 1364 1362 1139 925 941 928 926 ON31JI3VX1 $T=394800 168000 1 0 $X=394370 $Y=162880
X9113 1364 1362 266 278 284 788 EO3JI3VX1 $T=167440 141120 0 0 $X=167010 $Y=140480
X9114 1364 1362 266 279 289 1331 EO3JI3VX1 $T=169680 150080 1 0 $X=169250 $Y=144960
X9115 1364 1362 152 72 BUJI3VX2 $T=124880 194880 1 0 $X=124450 $Y=189760
X9116 1364 1362 312 350 BUJI3VX2 $T=192640 212800 0 0 $X=192210 $Y=212160
X9117 1364 1362 384 148 BUJI3VX2 $T=216160 33600 0 0 $X=215730 $Y=32960
X9118 1364 1362 367 152 BUJI3VX2 $T=220640 185920 1 0 $X=220210 $Y=180800
X9119 1364 1362 426 245 BUJI3VX2 $T=241920 33600 1 180 $X=238130 $Y=32960
X9120 1364 1362 433 191 BUJI3VX2 $T=268800 212800 1 180 $X=265010 $Y=212160
X9121 1364 1362 467 1405 BUJI3VX2 $T=282240 132160 0 0 $X=281810 $Y=131520
X9122 1364 1362 483 497 BUJI3VX2 $T=305760 203840 0 0 $X=305330 $Y=203200
X9123 1364 1362 531 up_switches<16> BUJI3VX2 $T=328160 24640 1 0 $X=327730 $Y=19520
X9124 1364 1362 527 up_switches<17> BUJI3VX2 $T=332080 24640 1 0 $X=331650 $Y=19520
X9125 1364 1362 549 up_switches<18> BUJI3VX2 $T=335440 24640 1 0 $X=335010 $Y=19520
X9126 1364 1362 869 up_switches<19> BUJI3VX2 $T=342720 24640 1 0 $X=342290 $Y=19520
X9127 1364 1362 876 up_switches<21> BUJI3VX2 $T=352240 24640 1 180 $X=348450 $Y=24000
X9128 1364 1362 579 up_switches<20> BUJI3VX2 $T=362880 24640 0 180 $X=359090 $Y=19520
X9129 1364 1362 577 up_switches<23> BUJI3VX2 $T=360640 33600 1 0 $X=360210 $Y=28480
X9130 1364 1362 908 up_switches<26> BUJI3VX2 $T=362880 24640 1 0 $X=362450 $Y=19520
X9131 1364 1362 898 up_switches<25> BUJI3VX2 $T=366800 24640 0 0 $X=366370 $Y=24000
X9132 1364 1362 887 up_switches<24> BUJI3VX2 $T=366800 33600 1 0 $X=366370 $Y=28480
X9133 1364 1362 1126 up_switches<27> BUJI3VX2 $T=370160 24640 0 0 $X=369730 $Y=24000
X9134 1364 1362 395 22 BUJI3VX2 $T=372960 51520 0 0 $X=372530 $Y=50880
X9135 1364 1362 603 up_switches<28> BUJI3VX2 $T=381360 24640 1 0 $X=380930 $Y=19520
X9136 1364 1362 597 up_switches<29> BUJI3VX2 $T=397600 24640 0 180 $X=393810 $Y=19520
X9137 1364 1362 1140 up_switches<30> BUJI3VX2 $T=402640 24640 0 180 $X=398850 $Y=19520
X9138 1364 1362 643 up_switches<31> BUJI3VX2 $T=402640 24640 1 0 $X=402210 $Y=19520
X9139 1364 1362 140 enable INJI3VX3 $T=92960 176960 0 0 $X=92530 $Y=176320
X9140 1364 1362 1026 165 INJI3VX3 $T=181440 159040 0 0 $X=181010 $Y=158400
X9141 1364 1362 245 662 INJI3VX3 $T=194880 33600 1 0 $X=194450 $Y=28480
X9142 1364 1362 1409 852 INJI3VX3 $T=215600 212800 0 0 $X=215170 $Y=212160
X9143 1364 1362 1061 378 INJI3VX3 $T=233520 159040 1 180 $X=230290 $Y=158400
X9144 1364 1362 488 up_switches<14> INJI3VX3 $T=303520 24640 1 0 $X=303090 $Y=19520
X9145 1364 1362 491 up_switches<15> INJI3VX3 $T=308560 24640 1 0 $X=308130 $Y=19520
X9146 1364 1362 938 up_switches<22> INJI3VX3 $T=325920 24640 0 0 $X=325490 $Y=24000
X9147 1364 1362 820 140 1087 1229 NA3I2JI3VX1 $T=216160 168000 1 180 $X=211810 $Y=167360
X9148 1364 1362 13 1057 824 1334 NA3I2JI3VX1 $T=220640 194880 0 180 $X=216290 $Y=189760
X9149 1364 1362 499 502 498 493 NA3I2JI3VX1 $T=311920 212800 1 180 $X=307570 $Y=212160
X9150 1364 1362 547 543 529 1410 NA3I2JI3VX1 $T=334880 168000 1 180 $X=330530 $Y=167360
X9151 1364 1362 304 279 1015 783 EN3JI3VX1 $T=183120 123200 1 180 $X=172050 $Y=122560
X9152 1364 1362 32 694 72 102 26 694 SDFRRQJI3VX1 $T=62160 78400 1 180 $X=41570 $Y=77760
X9153 1364 1362 28 84 72 128 26 84 SDFRRQJI3VX1 $T=62160 96320 0 180 $X=41570 $Y=91200
X9154 1364 1362 30 73 72 175 26 73 SDFRRQJI3VX1 $T=62160 96320 1 180 $X=41570 $Y=95680
X9155 1364 1362 32 108 72 126 26 108 SDFRRQJI3VX1 $T=62720 69440 1 180 $X=42130 $Y=68800
X9156 1364 1362 28 109 72 126 26 109 SDFRRQJI3VX1 $T=62720 78400 0 180 $X=42130 $Y=73280
X9157 1364 1362 28 695 72 102 26 695 SDFRRQJI3VX1 $T=62720 87360 0 180 $X=42130 $Y=82240
X9158 1364 1362 30 82 72 123 26 82 SDFRRQJI3VX1 $T=62720 105280 0 180 $X=42130 $Y=100160
X9159 1364 1362 30 110 72 103 26 110 SDFRRQJI3VX1 $T=62720 105280 1 180 $X=42130 $Y=104640
X9160 1364 1362 30 112 72 173 26 112 SDFRRQJI3VX1 $T=63280 114240 0 180 $X=42690 $Y=109120
X9161 1364 1362 30 95 72 127 26 95 SDFRRQJI3VX1 $T=77280 123200 1 180 $X=56690 $Y=122560
X9162 1364 1362 30 99 72 177 26 99 SDFRRQJI3VX1 $T=80080 123200 0 180 $X=59490 $Y=118080
X9163 1364 1362 30 107 72 126 26 107 SDFRRQJI3VX1 $T=80080 132160 0 180 $X=59490 $Y=127040
X9164 1364 1362 32 29 98 127 26 29 SDFRRQJI3VX1 $T=64960 78400 0 0 $X=64530 $Y=77760
X9165 1364 1362 28 958 72 127 26 958 SDFRRQJI3VX1 $T=64960 87360 1 0 $X=64530 $Y=82240
X9166 1364 1362 32 144 72 128 26 144 SDFRRQJI3VX1 $T=64960 87360 0 0 $X=64530 $Y=86720
X9167 1364 1362 26 103 72 123 33 103 SDFRRQJI3VX1 $T=65520 96320 1 0 $X=65090 $Y=91200
X9168 1364 1362 26 123 72 127 33 123 SDFRRQJI3VX1 $T=65520 96320 0 0 $X=65090 $Y=95680
X9169 1364 1362 26 127 72 126 33 127 SDFRRQJI3VX1 $T=65520 105280 0 0 $X=65090 $Y=104640
X9170 1364 1362 26 126 72 102 33 126 SDFRRQJI3VX1 $T=66080 105280 1 0 $X=65650 $Y=100160
X9171 1364 1362 26 102 72 128 33 102 SDFRRQJI3VX1 $T=67760 114240 0 0 $X=67330 $Y=113600
X9172 1364 1362 30 151 72 128 26 151 SDFRRQJI3VX1 $T=70560 159040 1 0 $X=70130 $Y=153920
X9173 1364 1362 30 716 72 102 26 716 SDFRRQJI3VX1 $T=71120 150080 0 0 $X=70690 $Y=149440
X9174 1364 1362 28 154 98 123 26 154 SDFRRQJI3VX1 $T=95200 69440 0 180 $X=74610 $Y=64320
X9175 1364 1362 32 718 98 123 26 718 SDFRRQJI3VX1 $T=95200 69440 1 180 $X=74610 $Y=68800
X9176 1364 1362 32 136 98 103 26 136 SDFRRQJI3VX1 $T=95200 78400 0 180 $X=74610 $Y=73280
X9177 1364 1362 659 127 72 137 26 137 SDFRRQJI3VX1 $T=95200 114240 0 180 $X=74610 $Y=109120
X9178 1364 1362 30 935 72 172 26 935 SDFRRQJI3VX1 $T=95200 132160 1 180 $X=74610 $Y=131520
X9179 1364 1362 659 126 72 719 26 719 SDFRRQJI3VX1 $T=95200 159040 1 180 $X=74610 $Y=158400
X9180 1364 1362 26 175 72 103 33 175 SDFRRQJI3VX1 $T=103040 69440 1 0 $X=102610 $Y=64320
X9181 1364 1362 28 969 98 103 26 969 SDFRRQJI3VX1 $T=103040 78400 1 0 $X=102610 $Y=73280
X9182 1364 1362 659 123 98 186 26 186 SDFRRQJI3VX1 $T=103040 105280 1 0 $X=102610 $Y=100160
X9183 1364 1362 26 128 72 160 33 128 SDFRRQJI3VX1 $T=103040 123200 0 0 $X=102610 $Y=122560
X9184 1364 1362 659 103 98 1188 26 1188 SDFRRQJI3VX1 $T=103040 132160 1 0 $X=102610 $Y=127040
X9185 1364 1362 30 1183 98 261 26 1183 SDFRRQJI3VX1 $T=103040 141120 0 0 $X=102610 $Y=140480
X9186 1364 1362 30 159 72 160 26 159 SDFRRQJI3VX1 $T=103040 159040 1 0 $X=102610 $Y=153920
X9187 1364 1362 659 102 406 161 SPI_CS 161 SDFRRQJI3VX1 $T=103040 185920 1 0 $X=102610 $Y=180800
X9188 1364 1362 659 128 72 162 SPI_CS 162 SDFRRQJI3VX1 $T=103040 185920 0 0 $X=102610 $Y=185280
X9189 1364 1362 659 175 98 200 26 200 SDFRRQJI3VX1 $T=110320 105280 0 0 $X=109890 $Y=104640
X9190 1364 1362 32 202 165 175 26 202 SDFRRQJI3VX1 $T=110880 69440 0 0 $X=110450 $Y=68800
X9191 1364 1362 32 171 165 173 26 171 SDFRRQJI3VX1 $T=110880 87360 1 0 $X=110450 $Y=82240
X9192 1364 1362 28 203 165 173 26 203 SDFRRQJI3VX1 $T=110880 87360 0 0 $X=110450 $Y=86720
X9193 1364 1362 26 172 165 177 33 172 SDFRRQJI3VX1 $T=110880 96320 1 0 $X=110450 $Y=91200
X9194 1364 1362 28 1189 98 175 26 1189 SDFRRQJI3VX1 $T=111440 78400 0 0 $X=111010 $Y=77760
X9195 1364 1362 659 177 98 182 26 182 SDFRRQJI3VX1 $T=113680 114240 1 0 $X=113250 $Y=109120
X9196 1364 1362 659 160 406 184 SPI_CS 184 SDFRRQJI3VX1 $T=115360 212800 0 0 $X=114930 $Y=212160
X9197 1364 1362 26 173 98 175 33 173 SDFRRQJI3VX1 $T=123200 96320 0 0 $X=122770 $Y=95680
X9198 1364 1362 659 173 98 750 26 750 SDFRRQJI3VX1 $T=123200 123200 0 0 $X=122770 $Y=122560
X9199 1364 1362 28 983 165 177 26 983 SDFRRQJI3VX1 $T=131600 78400 1 0 $X=131170 $Y=73280
X9200 1364 1362 32 209 165 177 26 209 SDFRRQJI3VX1 $T=131600 87360 1 0 $X=131170 $Y=82240
X9201 1364 1362 26 177 98 173 33 177 SDFRRQJI3VX1 $T=132160 105280 0 0 $X=131730 $Y=104640
X9202 1364 1362 32 1305 165 160 26 1305 SDFRRQJI3VX1 $T=142240 96320 1 0 $X=141810 $Y=91200
X9203 1364 1362 28 1013 165 172 26 1013 SDFRRQJI3VX1 $T=142800 78400 0 0 $X=142370 $Y=77760
X9204 1364 1362 28 238 165 160 26 238 SDFRRQJI3VX1 $T=142800 87360 0 0 $X=142370 $Y=86720
X9205 1364 1362 272 237 152 240 15 272 SDFRRQJI3VX1 $T=149520 176960 1 0 $X=149090 $Y=171840
X9206 1364 1362 1019 43 152 246 15 1019 SDFRRQJI3VX1 $T=152880 194880 0 0 $X=152450 $Y=194240
X9207 1364 1362 32 254 165 261 26 254 SDFRRQJI3VX1 $T=162400 78400 1 0 $X=161970 $Y=73280
X9208 1364 1362 32 255 165 172 26 255 SDFRRQJI3VX1 $T=162400 87360 1 0 $X=161970 $Y=82240
X9209 1364 1362 28 792 165 261 26 792 SDFRRQJI3VX1 $T=162960 69440 0 0 $X=162530 $Y=68800
X9210 1364 1362 26 261 165 172 33 261 SDFRRQJI3VX1 $T=165760 87360 0 0 $X=165330 $Y=86720
X9211 1364 1362 30 780 165 301 26 780 SDFRRQJI3VX1 $T=186480 96320 0 180 $X=165890 $Y=91200
X9212 1364 1362 32 789 165 301 26 789 SDFRRQJI3VX1 $T=178640 60480 0 0 $X=178210 $Y=59840
X9213 1364 1362 28 297 165 301 26 297 SDFRRQJI3VX1 $T=179760 69440 1 0 $X=179330 $Y=64320
X9214 1364 1362 32 1038 406 303 26 1038 SDFRRQJI3VX1 $T=183120 78400 1 0 $X=182690 $Y=73280
X9215 1364 1362 28 302 406 805 26 302 SDFRRQJI3VX1 $T=203280 78400 1 180 $X=182690 $Y=77760
X9216 1364 1362 26 303 152 301 33 303 SDFRRQJI3VX1 $T=183120 96320 0 0 $X=182690 $Y=95680
X9217 1364 1362 26 301 152 261 33 301 SDFRRQJI3VX1 $T=187040 87360 1 0 $X=186610 $Y=82240
X9218 1364 1362 28 309 406 303 41 309 SDFRRQJI3VX1 $T=188160 69440 0 0 $X=187730 $Y=68800
X9219 1364 1362 659 301 406 811 SPI_CS 811 SDFRRQJI3VX1 $T=212240 141120 0 180 $X=191650 $Y=136000
X9220 1364 1362 659 172 406 321 SPI_CS 321 SDFRRQJI3VX1 $T=193200 141120 0 0 $X=192770 $Y=140480
X9221 1364 1362 659 261 406 322 SPI_CS 322 SDFRRQJI3VX1 $T=193200 159040 0 0 $X=192770 $Y=158400
X9222 1364 1362 32 1056 406 363 41 1056 SDFRRQJI3VX1 $T=223440 78400 0 180 $X=202850 $Y=73280
X9223 1364 1362 32 366 406 805 41 366 SDFRRQJI3VX1 $T=223440 78400 1 180 $X=202850 $Y=77760
X9224 1364 1362 30 826 406 805 41 826 SDFRRQJI3VX1 $T=223440 87360 1 180 $X=202850 $Y=86720
X9225 1364 1362 41 363 152 805 33 363 SDFRRQJI3VX1 $T=223440 96320 0 180 $X=202850 $Y=91200
X9226 1364 1362 41 805 152 303 33 805 SDFRRQJI3VX1 $T=223440 96320 1 180 $X=202850 $Y=95680
X9227 1364 1362 30 325 406 303 41 325 SDFRRQJI3VX1 $T=223440 105280 0 180 $X=202850 $Y=100160
X9228 1364 1362 30 329 406 363 41 329 SDFRRQJI3VX1 $T=223440 105280 1 180 $X=202850 $Y=104640
X9229 1364 1362 30 337 406 376 41 337 SDFRRQJI3VX1 $T=223440 114240 0 180 $X=202850 $Y=109120
X9230 1364 1362 30 12 406 372 41 12 SDFRRQJI3VX1 $T=223440 123200 1 180 $X=202850 $Y=122560
X9231 1364 1362 659 303 406 823 41 823 SDFRRQJI3VX1 $T=223440 132160 0 180 $X=202850 $Y=127040
X9232 1364 1362 30 1232 406 469 41 1232 SDFRRQJI3VX1 $T=223440 132160 1 180 $X=202850 $Y=131520
X9233 1364 1362 28 828 378 363 41 828 SDFRRQJI3VX1 $T=231840 69440 0 0 $X=231410 $Y=68800
X9234 1364 1362 41 160 379 374 33 160 SDFRRQJI3VX1 $T=231840 212800 0 0 $X=231410 $Y=212160
X9235 1364 1362 32 829 378 372 41 829 SDFRRQJI3VX1 $T=232960 78400 0 0 $X=232530 $Y=77760
X9236 1364 1362 28 371 378 376 41 371 SDFRRQJI3VX1 $T=232960 87360 1 0 $X=232530 $Y=82240
X9237 1364 1362 28 830 378 372 41 830 SDFRRQJI3VX1 $T=232960 87360 0 0 $X=232530 $Y=86720
X9238 1364 1362 41 376 378 363 33 376 SDFRRQJI3VX1 $T=232960 96320 0 0 $X=232530 $Y=95680
X9239 1364 1362 659 805 395 375 41 375 SDFRRQJI3VX1 $T=232960 105280 0 0 $X=232530 $Y=104640
X9240 1364 1362 41 372 395 376 33 372 SDFRRQJI3VX1 $T=233520 105280 1 0 $X=233090 $Y=100160
X9241 1364 1362 659 363 395 382 41 382 SDFRRQJI3VX1 $T=237440 114240 0 0 $X=237010 $Y=113600
X9242 1364 1362 659 372 395 386 41 386 SDFRRQJI3VX1 $T=239680 123200 1 0 $X=239250 $Y=118080
X9243 1364 1362 28 427 378 415 41 427 SDFRRQJI3VX1 $T=267680 78400 0 180 $X=247090 $Y=73280
X9244 1364 1362 30 1086 406 415 SPI_CS 1086 SDFRRQJI3VX1 $T=271040 141120 0 180 $X=250450 $Y=136000
X9245 1364 1362 30 392 379 455 SPI_CS 392 SDFRRQJI3VX1 $T=271040 141120 1 180 $X=250450 $Y=140480
X9246 1364 1362 30 403 395 468 SPI_CS 403 SDFRRQJI3VX1 $T=272160 132160 1 180 $X=251570 $Y=131520
X9247 1364 1362 32 1078 378 376 41 1078 SDFRRQJI3VX1 $T=254800 87360 1 0 $X=254370 $Y=82240
X9248 1364 1362 28 847 378 469 41 847 SDFRRQJI3VX1 $T=254800 87360 0 0 $X=254370 $Y=86720
X9249 1364 1362 32 450 378 469 41 450 SDFRRQJI3VX1 $T=255360 96320 1 0 $X=254930 $Y=91200
X9250 1364 1362 659 376 395 451 41 451 SDFRRQJI3VX1 $T=255920 114240 1 0 $X=255490 $Y=109120
X9251 1364 1362 41 415 378 372 33 415 SDFRRQJI3VX1 $T=256480 105280 1 0 $X=256050 $Y=100160
X9252 1364 1362 32 444 378 415 41 444 SDFRRQJI3VX1 $T=271600 78400 1 0 $X=271170 $Y=73280
X9253 1364 1362 41 455 378 415 33 455 SDFRRQJI3VX1 $T=274400 96320 0 0 $X=273970 $Y=95680
X9254 1364 1362 32 1260 378 455 41 1260 SDFRRQJI3VX1 $T=274960 78400 0 0 $X=274530 $Y=77760
X9255 1364 1362 28 454 378 455 SPI_CS 454 SDFRRQJI3VX1 $T=274960 87360 1 0 $X=274530 $Y=82240
X9256 1364 1362 41 469 378 455 33 469 SDFRRQJI3VX1 $T=295120 87360 1 180 $X=274530 $Y=86720
X9257 1364 1362 659 469 395 863 SPI_CS 863 SDFRRQJI3VX1 $T=274960 132160 1 0 $X=274530 $Y=127040
X9258 1364 1362 659 415 395 461 SPI_CS 461 SDFRRQJI3VX1 $T=274960 141120 1 0 $X=274530 $Y=136000
X9259 1364 1362 659 455 395 481 SPI_CS 481 SDFRRQJI3VX1 $T=274960 141120 0 0 $X=274530 $Y=140480
X9260 1364 1362 30 443 395 466 SPI_CS 443 SDFRRQJI3VX1 $T=295120 150080 0 180 $X=274530 $Y=144960
X9261 1364 1362 41 460 379 463 33 460 SDFRRQJI3VX1 $T=275520 212800 1 0 $X=275090 $Y=207680
X9262 1364 1362 41 466 378 468 33 466 SDFRRQJI3VX1 $T=278880 105280 0 0 $X=278450 $Y=104640
X9263 1364 1362 41 468 378 469 33 468 SDFRRQJI3VX1 $T=278880 114240 1 0 $X=278450 $Y=109120
X9264 1364 1362 41 463 379 483 33 463 SDFRRQJI3VX1 $T=299040 203840 1 180 $X=278450 $Y=203200
X9265 1364 1362 1096 877 379 530 15 1096 SDFRRQJI3VX1 $T=310800 185920 0 180 $X=290210 $Y=180800
X9266 1364 1362 41 478 395 480 33 478 SDFRRQJI3VX1 $T=291760 168000 0 0 $X=291330 $Y=167360
X9267 1364 1362 41 479 395 478 33 472 SDFRRQJI3VX1 $T=291760 185920 0 0 $X=291330 $Y=185280
X9268 1364 1362 41 497 395 484 33 483 SDFRRQJI3VX1 $T=312480 203840 0 180 $X=291890 $Y=198720
X9269 1364 1362 32 501 378 468 41 501 SDFRRQJI3VX1 $T=292880 105280 1 0 $X=292450 $Y=100160
X9270 1364 1362 41 871 395 472 33 484 SDFRRQJI3VX1 $T=292880 194880 0 0 $X=292450 $Y=194240
X9271 1364 1362 41 480 395 496 33 480 SDFRRQJI3VX1 $T=314160 114240 1 180 $X=293570 $Y=113600
X9272 1364 1362 28 1100 378 468 41 1100 SDFRRQJI3VX1 $T=294560 96320 1 0 $X=294130 $Y=91200
X9273 1364 1362 28 505 378 466 41 505 SDFRRQJI3VX1 $T=295120 87360 1 0 $X=294690 $Y=82240
X9274 1364 1362 32 506 378 466 41 506 SDFRRQJI3VX1 $T=295120 87360 0 0 $X=294690 $Y=86720
X9275 1364 1362 41 504 378 466 33 504 SDFRRQJI3VX1 $T=295120 123200 1 0 $X=294690 $Y=118080
X9276 1364 1362 659 504 395 515 SPI_CS 515 SDFRRQJI3VX1 $T=298480 132160 1 0 $X=298050 $Y=127040
X9277 1364 1362 659 468 395 516 SPI_CS 516 SDFRRQJI3VX1 $T=298480 141120 1 0 $X=298050 $Y=136000
X9278 1364 1362 30 508 395 504 SPI_CS 508 SDFRRQJI3VX1 $T=318640 141120 1 180 $X=298050 $Y=140480
X9279 1364 1362 659 466 395 517 SPI_CS 517 SDFRRQJI3VX1 $T=298480 150080 1 0 $X=298050 $Y=144960
X9280 1364 1362 41 496 395 614 33 496 SDFRRQJI3VX1 $T=333760 114240 0 180 $X=313170 $Y=109120
X9281 1364 1362 32 546 395 504 SPI_CS 546 SDFRRQJI3VX1 $T=314720 96320 0 0 $X=314290 $Y=95680
X9282 1364 1362 41 511 395 504 33 511 SDFRRQJI3VX1 $T=314720 105280 1 0 $X=314290 $Y=100160
X9283 1364 1362 28 514 395 504 SPI_CS 514 SDFRRQJI3VX1 $T=315840 96320 1 0 $X=315410 $Y=91200
X9284 1364 1362 30 883 395 511 SPI_CS 883 SDFRRQJI3VX1 $T=316960 114240 0 0 $X=316530 $Y=113600
X9285 1364 1362 32 550 395 511 SPI_CS 550 SDFRRQJI3VX1 $T=338240 87360 0 180 $X=317650 $Y=82240
X9286 1364 1362 28 551 395 511 SPI_CS 551 SDFRRQJI3VX1 $T=338800 78400 1 180 $X=318210 $Y=77760
X9287 1364 1362 28 573 395 570 SPI_CS 573 SDFRRQJI3VX1 $T=351680 69440 1 180 $X=331090 $Y=68800
X9288 1364 1362 32 574 395 570 SPI_CS 574 SDFRRQJI3VX1 $T=351680 78400 0 180 $X=331090 $Y=73280
X9289 1364 1362 41 570 395 511 33 570 SDFRRQJI3VX1 $T=352240 87360 1 180 $X=331650 $Y=86720
X9290 1364 1362 30 541 395 584 SPI_CS 541 SDFRRQJI3VX1 $T=352240 105280 1 180 $X=331650 $Y=104640
X9291 1364 1362 30 1279 395 570 SPI_CS 1279 SDFRRQJI3VX1 $T=352240 123200 0 180 $X=331650 $Y=118080
X9292 1364 1362 30 20 395 583 SPI_CS 20 SDFRRQJI3VX1 $T=352240 123200 1 180 $X=331650 $Y=122560
X9293 1364 1362 32 1136 22 583 SPI_CS 1136 SDFRRQJI3VX1 $T=360080 69440 0 0 $X=359650 $Y=68800
X9294 1364 1362 28 600 22 583 SPI_CS 600 SDFRRQJI3VX1 $T=360080 78400 1 0 $X=359650 $Y=73280
X9295 1364 1362 32 907 22 584 SPI_CS 907 SDFRRQJI3VX1 $T=360080 78400 0 0 $X=359650 $Y=77760
X9296 1364 1362 28 580 22 584 SPI_CS 580 SDFRRQJI3VX1 $T=360080 87360 1 0 $X=359650 $Y=82240
X9297 1364 1362 41 584 22 570 33 584 SDFRRQJI3VX1 $T=360080 87360 0 0 $X=359650 $Y=86720
X9298 1364 1362 41 585 22 583 33 585 SDFRRQJI3VX1 $T=360080 96320 1 0 $X=359650 $Y=91200
X9299 1364 1362 41 583 22 584 33 583 SDFRRQJI3VX1 $T=360080 96320 0 0 $X=359650 $Y=95680
X9300 1364 1362 30 601 22 582 SPI_CS 601 SDFRRQJI3VX1 $T=360080 114240 0 0 $X=359650 $Y=113600
X9301 1364 1362 30 602 22 585 SPI_CS 602 SDFRRQJI3VX1 $T=360080 123200 1 0 $X=359650 $Y=118080
X9302 1364 1362 30 1293 22 578 SPI_CS 1293 SDFRRQJI3VX1 $T=360080 123200 0 0 $X=359650 $Y=122560
X9303 1364 1362 30 1137 22 614 SPI_CS 1137 SDFRRQJI3VX1 $T=360080 132160 1 0 $X=359650 $Y=127040
X9304 1364 1362 41 582 22 585 33 582 SDFRRQJI3VX1 $T=361200 105280 1 0 $X=360770 $Y=100160
X9305 1364 1362 41 578 22 582 33 578 SDFRRQJI3VX1 $T=381360 105280 1 180 $X=360770 $Y=104640
X9306 1364 1362 41 614 22 578 33 614 SDFRRQJI3VX1 $T=381360 114240 0 180 $X=360770 $Y=109120
X9307 1364 1362 28 917 22 614 SPI_CS 917 SDFRRQJI3VX1 $T=380240 78400 0 0 $X=379810 $Y=77760
X9308 1364 1362 32 681 22 614 SPI_CS 681 SDFRRQJI3VX1 $T=380240 87360 1 0 $X=379810 $Y=82240
X9309 1364 1362 32 682 22 585 SPI_CS 682 SDFRRQJI3VX1 $T=380240 87360 0 0 $X=379810 $Y=86720
X9310 1364 1362 28 611 22 585 SPI_CS 611 SDFRRQJI3VX1 $T=380240 96320 0 0 $X=379810 $Y=95680
X9311 1364 1362 642 634 22 633 19 633 SDFRRQJI3VX1 $T=391440 132160 0 0 $X=391010 $Y=131520
X9312 1364 1362 32 23 22 578 SPI_CS 23 SDFRRQJI3VX1 $T=395360 78400 1 0 $X=394930 $Y=73280
X9313 1364 1362 32 638 22 582 SPI_CS 638 SDFRRQJI3VX1 $T=395360 96320 1 0 $X=394930 $Y=91200
X9314 1364 1362 28 1150 22 578 SPI_CS 1150 SDFRRQJI3VX1 $T=400400 87360 1 0 $X=399970 $Y=82240
X9315 1364 1362 28 24 22 582 SPI_CS 24 SDFRRQJI3VX1 $T=400400 87360 0 0 $X=399970 $Y=86720
X9316 1364 1362 946 1154 79 NO2JI3VX0 $T=40880 168000 1 180 $X=38210 $Y=167360
X9317 1364 1362 945 131 697 NO2JI3VX0 $T=44800 159040 0 0 $X=44370 $Y=158400
X9318 1364 1362 69 94 699 NO2JI3VX0 $T=47040 159040 1 0 $X=46610 $Y=153920
X9319 1364 1362 951 93 692 NO2JI3VX0 $T=53200 168000 1 180 $X=50530 $Y=167360
X9320 1364 1362 653 952 1165 NO2JI3VX0 $T=52640 176960 0 0 $X=52210 $Y=176320
X9321 1364 1362 93 97 952 NO2JI3VX0 $T=53760 168000 1 0 $X=53330 $Y=162880
X9322 1364 1362 118 1169 111 NO2JI3VX0 $T=62720 185920 0 180 $X=60050 $Y=180800
X9323 1364 1362 85 711 120 NO2JI3VX0 $T=62160 159040 1 0 $X=61730 $Y=153920
X9324 1364 1362 129 714 135 NO2JI3VX0 $T=69440 185920 0 180 $X=66770 $Y=180800
X9325 1364 1362 129 960 122 NO2JI3VX0 $T=71680 203840 0 180 $X=69010 $Y=198720
X9326 1364 1362 96 1178 132 NO2JI3VX0 $T=77840 194880 1 0 $X=77410 $Y=189760
X9327 1364 1362 1178 139 140 NO2JI3VX0 $T=80640 185920 1 180 $X=77970 $Y=185280
X9328 1364 1362 761 1002 776 NO2JI3VX0 $T=148960 123200 1 0 $X=148530 $Y=118080
X9329 1364 1362 272 1377 1022 NO2JI3VX0 $T=179200 176960 1 180 $X=176530 $Y=176320
X9330 1364 1362 793 310 292 NO2JI3VX0 $T=179760 203840 1 0 $X=179330 $Y=198720
X9331 1364 1362 1411 1029 40 NO2JI3VX0 $T=184800 185920 1 0 $X=184370 $Y=180800
X9332 1364 1362 790 333 807 NO2JI3VX0 $T=204960 185920 1 180 $X=202290 $Y=185280
X9333 1364 1362 51 1392 810 NO2JI3VX0 $T=218960 176960 0 180 $X=216290 $Y=171840
X9334 1364 1362 666 356 14 NO2JI3VX0 $T=220080 185920 0 180 $X=217410 $Y=180800
X9335 1364 1362 834 1068 383 NO2JI3VX0 $T=239680 168000 1 0 $X=239250 $Y=162880
X9336 1364 1362 53 1070 1239 NO2JI3VX0 $T=240240 194880 0 0 $X=239810 $Y=194240
X9337 1364 1362 423 53 377 NO2JI3VX0 $T=244720 194880 1 180 $X=242050 $Y=194240
X9338 1364 1362 1063 841 834 NO2JI3VX0 $T=245280 176960 0 180 $X=242610 $Y=171840
X9339 1364 1362 844 404 397 NO2JI3VX0 $T=253120 176960 1 180 $X=250450 $Y=176320
X9340 1364 1362 1241 401 844 NO2JI3VX0 $T=253120 185920 0 180 $X=250450 $Y=180800
X9341 1364 1362 410 1080 846 NO2JI3VX0 $T=255360 168000 0 0 $X=254930 $Y=167360
X9342 1364 1362 1082 416 414 NO2JI3VX0 $T=261520 185920 0 180 $X=258850 $Y=180800
X9343 1364 1362 527 886 531 NO2JI3VX0 $T=324800 24640 1 0 $X=324370 $Y=19520
X9344 1364 1362 1410 1343 1282 NO2JI3VX0 $T=330960 168000 1 180 $X=328290 $Y=167360
X9345 1364 1362 556 892 561 NO2JI3VX0 $T=337680 159040 1 0 $X=337250 $Y=153920
X9346 1364 1362 869 558 549 NO2JI3VX0 $T=338800 24640 0 0 $X=338370 $Y=24000
X9347 1364 1362 1402 1345 557 NO2JI3VX0 $T=339360 212800 0 0 $X=338930 $Y=212160
X9348 1364 1362 900 899 556 NO2JI3VX0 $T=343840 176960 1 180 $X=341170 $Y=176320
X9349 1364 1362 566 557 1389 NO2JI3VX0 $T=349440 212800 1 180 $X=346770 $Y=212160
X9350 1364 1362 571 1158 905 NO2JI3VX0 $T=352240 159040 1 180 $X=349570 $Y=158400
X9351 1364 1362 597 59 603 NO2JI3VX0 $T=380240 24640 0 180 $X=377570 $Y=19520
X9352 1364 1362 617 1386 626 NO2JI3VX0 $T=384720 114240 0 0 $X=384290 $Y=113600
X9353 1364 1362 624 1365 619 NO2JI3VX0 $T=384720 141120 0 0 $X=384290 $Y=140480
X9354 1364 1362 616 1352 553 NO2JI3VX0 $T=385280 159040 1 0 $X=384850 $Y=153920
X9355 1364 1362 620 617 633 NO2JI3VX0 $T=392000 105280 1 180 $X=389330 $Y=104640
X9356 1364 1362 643 904 1140 NO2JI3VX0 $T=393680 24640 0 180 $X=391010 $Y=19520
X9357 1364 1362 2 27 702 956 1163 NA4JI3VX0 $T=54320 159040 1 180 $X=49970 $Y=158400
X9358 1364 1362 1412 806 324 332 804 NA4JI3VX0 $T=198240 185920 1 0 $X=197810 $Y=180800
X9359 1364 1362 904 565 558 886 59 NA4JI3VX0 $T=347760 24640 1 0 $X=347330 $Y=19520
X9360 1364 1362 1141 1413 627 622 625 NA4JI3VX0 $T=394240 141120 0 180 $X=389890 $Y=136000
X9361 1364 1362 75 1414 68 NA2JI3VX0 $T=26320 168000 1 0 $X=25890 $Y=162880
X9362 1364 1362 83 1406 1159 NA2JI3VX0 $T=33600 150080 0 0 $X=33170 $Y=149440
X9363 1364 1362 75 1407 87 NA2JI3VX0 $T=42000 176960 1 180 $X=39330 $Y=176320
X9364 1364 1362 693 949 948 NA2JI3VX0 $T=40880 159040 0 0 $X=40450 $Y=158400
X9365 1364 1362 1369 86 1160 NA2JI3VX0 $T=42000 150080 0 0 $X=41570 $Y=149440
X9366 1364 1362 699 702 69 NA2JI3VX0 $T=49840 150080 1 180 $X=47170 $Y=149440
X9367 1364 1362 697 956 945 NA2JI3VX0 $T=47600 159040 0 0 $X=47170 $Y=158400
X9368 1364 1362 700 652 1169 NA2JI3VX0 $T=52080 185920 1 0 $X=51650 $Y=180800
X9369 1364 1362 952 705 92 NA2JI3VX0 $T=53760 176960 1 0 $X=53330 $Y=171840
X9370 1364 1362 120 713 85 NA2JI3VX0 $T=67760 159040 0 180 $X=65090 $Y=153920
X9371 1364 1362 1394 959 1171 NA2JI3VX0 $T=71120 168000 1 180 $X=68450 $Y=167360
X9372 1364 1362 157 147 148 NA2JI3VX0 $T=90160 24640 1 180 $X=87490 $Y=24000
X9373 1364 1362 721 1329 148 NA2JI3VX0 $T=91280 42560 0 180 $X=88610 $Y=37440
X9374 1364 1362 153 149 148 NA2JI3VX0 $T=92400 42560 1 0 $X=91970 $Y=37440
X9375 1364 1362 724 734 148 NA2JI3VX0 $T=103600 24640 0 0 $X=103170 $Y=24000
X9376 1364 1362 164 737 148 NA2JI3VX0 $T=110320 24640 1 180 $X=107650 $Y=24000
X9377 1364 1362 174 746 148 NA2JI3VX0 $T=115360 24640 1 180 $X=112690 $Y=24000
X9378 1364 1362 192 1190 148 NA2JI3VX0 $T=124880 33600 1 0 $X=124450 $Y=28480
X9379 1364 1362 205 756 148 NA2JI3VX0 $T=135520 33600 1 180 $X=132850 $Y=32960
X9380 1364 1362 210 982 212 NA2JI3VX0 $T=133280 114240 0 0 $X=132850 $Y=113600
X9381 1364 1362 198 222 212 NA2JI3VX0 $T=143920 114240 0 0 $X=143490 $Y=113600
X9382 1364 1362 226 224 148 NA2JI3VX0 $T=147840 24640 1 180 $X=145170 $Y=24000
X9383 1364 1362 1201 7 492 NA2JI3VX0 $T=148400 114240 1 180 $X=145730 $Y=113600
X9384 1364 1362 1355 227 492 NA2JI3VX0 $T=148960 123200 0 180 $X=146290 $Y=118080
X9385 1364 1362 763 769 148 NA2JI3VX0 $T=148960 33600 0 0 $X=148530 $Y=32960
X9386 1364 1362 997 1001 212 NA2JI3VX0 $T=148960 114240 1 0 $X=148530 $Y=109120
X9387 1364 1362 989 38 212 NA2JI3VX0 $T=152320 105280 0 0 $X=151890 $Y=104640
X9388 1364 1362 252 1156 148 NA2JI3VX0 $T=160720 33600 0 180 $X=158050 $Y=28480
X9389 1364 1362 1011 1008 492 NA2JI3VX0 $T=161840 114240 0 180 $X=159170 $Y=109120
X9390 1364 1362 966 1308 212 NA2JI3VX0 $T=164640 114240 1 0 $X=164210 $Y=109120
X9391 1364 1362 271 1307 148 NA2JI3VX0 $T=170240 33600 1 0 $X=169810 $Y=28480
X9392 1364 1362 286 1213 212 NA2JI3VX0 $T=175840 123200 1 0 $X=175410 $Y=118080
X9393 1364 1362 295 290 293 NA2JI3VX0 $T=183680 194880 0 180 $X=181010 $Y=189760
X9394 1364 1362 296 294 148 NA2JI3VX0 $T=182560 33600 0 0 $X=182130 $Y=32960
X9395 1364 1362 790 1332 1415 NA2JI3VX0 $T=183120 176960 1 0 $X=182690 $Y=171840
X9396 1364 1362 340 797 1415 NA2JI3VX0 $T=189280 176960 0 180 $X=186610 $Y=171840
X9397 1364 1362 798 308 300 NA2JI3VX0 $T=189840 194880 1 180 $X=187170 $Y=194240
X9398 1364 1362 317 315 1379 NA2JI3VX0 $T=195440 176960 1 0 $X=195010 $Y=171840
X9399 1364 1362 807 1219 790 NA2JI3VX0 $T=202160 185920 1 180 $X=199490 $Y=185280
X9400 1364 1362 335 326 148 NA2JI3VX0 $T=203280 42560 1 180 $X=200610 $Y=41920
X9401 1364 1362 328 349 46 NA2JI3VX0 $T=206080 203840 0 0 $X=205650 $Y=203200
X9402 1364 1362 813 344 148 NA2JI3VX0 $T=211120 33600 1 180 $X=208450 $Y=32960
X9403 1364 1362 45 1416 360 NA2JI3VX0 $T=211120 185920 0 180 $X=208450 $Y=180800
X9404 1364 1362 reset_l 1409 816 NA2JI3VX0 $T=211680 212800 0 0 $X=211250 $Y=212160
X9405 1364 1362 1045 1231 1050 NA2JI3VX0 $T=212800 203840 1 0 $X=212370 $Y=198720
X9406 1364 1362 381 817 384 NA2JI3VX0 $T=213920 33600 0 0 $X=213490 $Y=32960
X9407 1364 1362 14 360 1392 NA2JI3VX0 $T=216720 176960 0 180 $X=214050 $Y=171840
X9408 1364 1362 45 347 356 NA2JI3VX0 $T=220080 159040 1 0 $X=219650 $Y=153920
X9409 1364 1362 1066 831 384 NA2JI3VX0 $T=235760 33600 0 180 $X=233090 $Y=28480
X9410 1364 1362 1060 1233 1050 NA2JI3VX0 $T=237440 203840 0 180 $X=234770 $Y=198720
X9411 1364 1362 832 1338 384 NA2JI3VX0 $T=244160 33600 0 180 $X=241490 $Y=28480
X9412 1364 1362 1073 840 385 NA2JI3VX0 $T=248080 168000 1 180 $X=245410 $Y=167360
X9413 1364 1362 839 1241 841 NA2JI3VX0 $T=248640 185920 0 180 $X=245970 $Y=180800
X9414 1364 1362 399 1320 384 NA2JI3VX0 $T=253120 33600 0 0 $X=252690 $Y=32960
X9415 1364 1362 1066 848 462 NA2JI3VX0 $T=257040 42560 1 0 $X=256610 $Y=37440
X9416 1364 1362 413 1340 384 NA2JI3VX0 $T=261520 33600 1 0 $X=261090 $Y=28480
X9417 1364 1362 432 854 431 NA2JI3VX0 $T=269920 185920 1 180 $X=267250 $Y=185280
X9418 1364 1362 17 855 421 NA2JI3VX0 $T=268800 194880 1 0 $X=268370 $Y=189760
X9419 1364 1362 1381 858 856 NA2JI3VX0 $T=270480 176960 0 0 $X=270050 $Y=176320
X9420 1364 1362 441 859 384 NA2JI3VX0 $T=272160 42560 1 0 $X=271730 $Y=37440
X9421 1364 1362 456 452 449 NA2JI3VX0 $T=277760 185920 0 180 $X=275090 $Y=180800
X9422 1364 1362 447 862 449 NA2JI3VX0 $T=275520 185920 0 0 $X=275090 $Y=185280
X9423 1364 1362 457 440 384 NA2JI3VX0 $T=278320 33600 0 180 $X=275650 $Y=28480
X9424 1364 1362 458 853 384 NA2JI3VX0 $T=278320 42560 0 180 $X=275650 $Y=37440
X9425 1364 1362 453 865 384 NA2JI3VX0 $T=278320 24640 0 0 $X=277890 $Y=24000
X9426 1364 1362 45 1227 482 NA2JI3VX0 $T=281120 168000 0 0 $X=280690 $Y=167360
X9427 1364 1362 458 866 462 NA2JI3VX0 $T=282240 42560 1 0 $X=281810 $Y=37440
X9428 1364 1362 457 470 462 NA2JI3VX0 $T=282800 33600 1 0 $X=282370 $Y=28480
X9429 1364 1362 474 1264 384 NA2JI3VX0 $T=295680 24640 1 180 $X=293010 $Y=24000
X9430 1364 1362 1098 1265 384 NA2JI3VX0 $T=295680 33600 1 180 $X=293010 $Y=32960
X9431 1364 1362 45 1417 487 NA2JI3VX0 $T=297920 176960 1 0 $X=297490 $Y=171840
X9432 1364 1362 496 486 485 NA2JI3VX0 $T=302960 123200 0 0 $X=302530 $Y=122560
X9433 1364 1362 513 879 384 NA2JI3VX0 $T=313040 33600 1 180 $X=310370 $Y=32960
X9434 1364 1362 502 489 509 NA2JI3VX0 $T=313040 212800 0 0 $X=312610 $Y=212160
X9435 1364 1362 503 882 384 NA2JI3VX0 $T=316960 33600 1 0 $X=316530 $Y=28480
X9436 1364 1362 528 525 884 NA2JI3VX0 $T=321440 168000 1 0 $X=321010 $Y=162880
X9437 1364 1362 534 545 1281 NA2JI3VX0 $T=329840 176960 0 0 $X=329410 $Y=176320
X9438 1364 1362 544 891 542 NA2JI3VX0 $T=330960 194880 1 0 $X=330530 $Y=189760
X9439 1364 1362 535 889 384 NA2JI3VX0 $T=332080 33600 0 0 $X=331650 $Y=32960
X9440 1364 1362 537 1287 384 NA2JI3VX0 $T=337120 33600 1 0 $X=336690 $Y=28480
X9441 1364 1362 535 56 462 NA2JI3VX0 $T=337120 42560 1 0 $X=336690 $Y=37440
X9442 1364 1362 560 1384 462 NA2JI3VX0 $T=343280 42560 1 0 $X=342850 $Y=37440
X9443 1364 1362 560 1291 384 NA2JI3VX0 $T=345520 42560 1 0 $X=345090 $Y=37440
X9444 1364 1362 1128 906 384 NA2JI3VX0 $T=349440 51520 1 0 $X=349010 $Y=46400
X9445 1364 1362 905 567 571 NA2JI3VX0 $T=351680 168000 0 180 $X=349010 $Y=162880
X9446 1364 1362 587 897 1123 NA2JI3VX0 $T=365680 176960 0 180 $X=363010 $Y=171840
X9447 1364 1362 581 586 588 NA2JI3VX0 $T=363440 185920 1 0 $X=363010 $Y=180800
X9448 1364 1362 909 60 588 NA2JI3VX0 $T=367920 185920 0 180 $X=365250 $Y=180800
X9449 1364 1362 678 1347 384 NA2JI3VX0 $T=366240 42560 1 0 $X=365810 $Y=37440
X9450 1364 1362 61 1348 384 NA2JI3VX0 $T=370720 42560 0 180 $X=368050 $Y=37440
X9451 1364 1362 678 1349 462 NA2JI3VX0 $T=372960 42560 0 180 $X=370290 $Y=37440
X9452 1364 1362 590 1131 384 NA2JI3VX0 $T=371840 33600 1 0 $X=371410 $Y=28480
X9453 1364 1362 598 1361 384 NA2JI3VX0 $T=375200 42560 0 180 $X=372530 $Y=37440
X9454 1364 1362 598 1135 462 NA2JI3VX0 $T=376880 42560 1 0 $X=376450 $Y=37440
X9455 1364 1362 595 1327 384 NA2JI3VX0 $T=377440 33600 0 0 $X=377010 $Y=32960
X9456 1364 1362 606 610 1385 NA2JI3VX0 $T=385840 159040 1 180 $X=383170 $Y=158400
X9457 1364 1362 626 1408 621 NA2JI3VX0 $T=385840 123200 1 0 $X=385410 $Y=118080
X9458 1364 1362 618 622 606 NA2JI3VX0 $T=389200 141120 0 180 $X=386530 $Y=136000
X9459 1364 1362 635 1143 384 NA2JI3VX0 $T=396480 33600 0 180 $X=393810 $Y=28480
X9460 1364 1362 637 921 384 NA2JI3VX0 $T=396480 33600 1 180 $X=393810 $Y=32960
X9461 1364 1362 607 627 925 NA2JI3VX0 $T=395360 150080 1 0 $X=394930 $Y=144960
X9462 1364 1362 1139 926 1146 NA2JI3VX0 $T=395920 159040 0 0 $X=395490 $Y=158400
X9463 1364 1362 1147 642 1413 NA2JI3VX0 $T=402080 141120 0 180 $X=399410 $Y=136000
X9464 1364 1362 1418 662 149 down_switches<4> ON21JI3VX4 $T=91280 42560 1 180 $X=82450 $Y=41920
X9465 1364 1362 31 662 147 down_switches<1> ON21JI3VX4 $T=84560 24640 1 0 $X=84130 $Y=19520
X9466 1364 1362 1419 662 1329 down_switches<2> ON21JI3VX4 $T=87360 33600 0 0 $X=86930 $Y=32960
X9467 1364 1362 968 662 734 down_switches<3> ON21JI3VX4 $T=109760 24640 0 180 $X=100930 $Y=19520
X9468 1364 1362 736 662 737 down_switches<5> ON21JI3VX4 $T=109760 24640 1 0 $X=109330 $Y=19520
X9469 1364 1362 743 662 746 down_switches<6> ON21JI3VX4 $T=118160 24640 1 0 $X=117730 $Y=19520
X9470 1364 1362 977 662 1190 down_switches<7> ON21JI3VX4 $T=134960 24640 0 180 $X=126130 $Y=19520
X9471 1364 1362 760 662 756 down_switches<9> ON21JI3VX4 $T=137200 33600 0 180 $X=128370 $Y=28480
X9472 1364 1362 1420 662 224 down_switches<8> ON21JI3VX4 $T=140000 24640 1 180 $X=131170 $Y=24000
X9473 1364 1362 241 662 769 down_switches<0> ON21JI3VX4 $T=154560 33600 0 180 $X=145730 $Y=28480
X9474 1364 1362 1421 662 1156 down_switches<10> ON21JI3VX4 $T=160720 24640 0 180 $X=151890 $Y=19520
X9475 1364 1362 270 662 1307 down_switches<11> ON21JI3VX4 $T=170240 24640 1 180 $X=161410 $Y=24000
X9476 1364 1362 1422 662 294 down_switches<12> ON21JI3VX4 $T=183120 33600 0 180 $X=174290 $Y=28480
X9477 1364 1362 345 662 326 down_switches<13> ON21JI3VX4 $T=201600 42560 0 180 $X=192770 $Y=37440
X9478 1364 1362 1042 662 344 down_switches<14> ON21JI3VX4 $T=207760 33600 0 180 $X=198930 $Y=28480
X9479 1364 1362 1423 662 817 down_switches<15> ON21JI3VX4 $T=218960 33600 0 180 $X=210130 $Y=28480
X9480 1364 1362 1316 662 831 down_switches<17> ON21JI3VX4 $T=239120 24640 0 180 $X=230290 $Y=19520
X9481 1364 1362 1424 662 1338 down_switches<16> ON21JI3VX4 $T=241360 24640 1 180 $X=232530 $Y=24000
X9482 1364 1362 1425 662 1340 down_switches<20> ON21JI3VX4 $T=266560 24640 1 180 $X=257730 $Y=24000
X9483 1364 1362 1089 662 853 down_switches<18> ON21JI3VX4 $T=270480 42560 0 180 $X=261650 $Y=37440
X9484 1364 1362 1426 662 440 down_switches<19> ON21JI3VX4 $T=274960 33600 1 180 $X=266130 $Y=32960
X9485 1364 1362 1427 662 1264 down_switches<21> ON21JI3VX4 $T=296240 24640 0 180 $X=287410 $Y=19520
X9486 1364 1362 1099 662 1265 down_switches<22> ON21JI3VX4 $T=296240 33600 0 180 $X=287410 $Y=28480
X9487 1364 1362 510 662 879 down_switches<23> ON21JI3VX4 $T=317520 24640 1 180 $X=308690 $Y=24000
X9488 1364 1362 1108 662 882 down_switches<24> ON21JI3VX4 $T=322000 24640 0 180 $X=313170 $Y=19520
X9489 1364 1362 890 662 889 down_switches<25> ON21JI3VX4 $T=337120 24640 1 180 $X=328290 $Y=24000
X9490 1364 1362 568 662 1291 down_switches<26> ON21JI3VX4 $T=351120 33600 1 180 $X=342290 $Y=32960
X9491 1364 1362 1428 662 1347 down_switches<27> ON21JI3VX4 $T=366240 33600 1 180 $X=357410 $Y=32960
X9492 1364 1362 1294 662 1361 down_switches<28> ON21JI3VX4 $T=366240 42560 0 180 $X=357410 $Y=37440
X9493 1364 1362 593 662 1131 down_switches<31> ON21JI3VX4 $T=376880 24640 0 180 $X=368050 $Y=19520
X9494 1364 1362 630 662 921 down_switches<30> ON21JI3VX4 $T=393680 33600 1 180 $X=384850 $Y=32960
X9495 1364 1362 1429 662 1143 down_switches<29> ON21JI3VX4 $T=386960 24640 0 0 $X=386530 $Y=24000
X9496 1364 1362 115 210 1366 AND2JI3VX1 $T=61600 33600 1 0 $X=61170 $Y=28480
X9497 1364 1362 115 198 125 AND2JI3VX1 $T=62160 24640 0 0 $X=61730 $Y=24000
X9498 1364 1362 115 966 1367 AND2JI3VX1 $T=75600 33600 1 0 $X=75170 $Y=28480
X9499 1364 1362 115 989 725 AND2JI3VX1 $T=137760 33600 1 0 $X=137330 $Y=28480
X9500 1364 1362 115 997 726 AND2JI3VX1 $T=142240 24640 0 0 $X=141810 $Y=24000
X9501 1364 1362 115 286 287 AND2JI3VX1 $T=180320 24640 1 180 $X=176530 $Y=24000
X9502 1364 1362 343 938 488 491 559 NA4JI3VX2 $T=306320 24640 1 180 $X=298610 $Y=24000
X9503 1364 1362 462 426 384 NO2I1JI3VX2 $T=313040 33600 0 180 $X=307570 $Y=28480
X9504 1364 1362 1002 1199 216 EO2JI3VX0 $T=141680 123200 0 180 $X=135650 $Y=118080
X9505 1364 1362 1391 239 1430 EO2JI3VX0 $T=156240 132160 0 180 $X=150210 $Y=127040
X9506 1364 1362 295 293 1403 EO2JI3VX0 $T=181440 194880 0 180 $X=175410 $Y=189760
X9507 1364 1362 328 46 1404 EO2JI3VX0 $T=194320 203840 0 0 $X=193890 $Y=203200
X9508 1364 1362 17 421 448 EO2JI3VX0 $T=271040 203840 1 0 $X=270610 $Y=198720
X9509 1364 1362 460 IC_addr<1> 477 EO2JI3VX0 $T=278880 212800 0 0 $X=278450 $Y=212160
X9510 1364 1362 463 IC_addr<0> 1398 EO2JI3VX0 $T=286720 212800 0 0 $X=286290 $Y=212160
X9511 1364 1362 534 1281 522 EO2JI3VX0 $T=328160 176960 0 180 $X=322130 $Y=171840
X9512 1364 1362 79 691 90 AND2JI3VX0 $T=41440 168000 0 0 $X=41010 $Y=167360
X9513 1364 1362 105 713 1163 AND2JI3VX0 $T=61600 159040 0 180 $X=57810 $Y=153920
X9514 1364 1362 47 1270 1230 AND2JI3VX0 $T=211680 168000 1 0 $X=211250 $Y=162880
X9515 1364 1362 844 397 389 AND2JI3VX0 $T=250320 176960 1 180 $X=246530 $Y=176320
X9516 1364 1362 401 393 1401 AND2JI3VX0 $T=250880 194880 0 0 $X=250450 $Y=194240
X9517 1364 1362 462 832 1244 AND2JI3VX0 $T=255920 33600 0 180 $X=252130 $Y=28480
X9518 1364 1362 566 676 1402 AND2JI3VX0 $T=346640 212800 1 180 $X=342850 $Y=212160
X9519 1364 1362 462 590 608 AND2JI3VX0 $T=384160 33600 0 180 $X=380370 $Y=28480
X9520 1364 1362 919 622 616 AND2JI3VX0 $T=389200 150080 0 180 $X=385410 $Y=144960
X9521 1364 1362 462 635 927 AND2JI3VX0 $T=397040 33600 1 0 $X=396610 $Y=28480
X9522 1364 1362 462 637 932 AND2JI3VX0 $T=400400 33600 0 0 $X=399970 $Y=32960
X9523 1364 1362 653 1169 1167 111 700 AN22JI3VX1 $T=59360 185920 0 180 $X=55010 $Y=180800
X9524 1364 1362 132 960 124 129 122 AN22JI3VX1 $T=71680 194880 1 180 $X=67330 $Y=194240
X9525 1364 1362 135 129 957 134 133 AN22JI3VX1 $T=74480 176960 1 180 $X=70130 $Y=176320
X9526 1364 1362 216 231 1375 353 979 AN22JI3VX1 $T=137200 114240 0 0 $X=136770 $Y=113600
X9527 1364 1362 1193 231 988 353 981 AN22JI3VX1 $T=142240 132160 0 180 $X=137890 $Y=127040
X9528 1364 1362 1430 231 37 353 223 AN22JI3VX1 $T=150080 132160 0 180 $X=145730 $Y=127040
X9529 1364 1362 298 492 1007 353 236 AN22JI3VX1 $T=154560 123200 1 0 $X=154130 $Y=118080
X9530 1364 1362 277 492 273 353 264 AN22JI3VX1 $T=172480 132160 0 180 $X=168130 $Y=127040
X9531 1364 1362 304 492 1025 353 278 AN22JI3VX1 $T=184240 132160 0 180 $X=179890 $Y=127040
X9532 1364 1362 299 795 1032 793 292 AN22JI3VX1 $T=187040 203840 0 180 $X=182690 $Y=198720
X9533 1364 1362 813 245 488 148 346 AN22JI3VX1 $T=223440 33600 1 180 $X=219090 $Y=32960
X9534 1364 1362 807 1045 824 50 390 AN22JI3VX1 $T=223440 185920 1 180 $X=219090 $Y=185280
X9535 1364 1362 381 245 491 384 364 AN22JI3VX1 $T=240800 33600 0 180 $X=236450 $Y=28480
X9536 1364 1362 383 834 405 1063 837 AN22JI3VX1 $T=238000 159040 0 0 $X=237570 $Y=158400
X9537 1364 1362 385 841 1317 834 839 AN22JI3VX1 $T=241920 176960 0 0 $X=241490 $Y=176320
X9538 1364 1362 410 401 400 393 844 AN22JI3VX1 $T=254240 185920 1 180 $X=249890 $Y=185280
X9539 1364 1362 1098 426 938 384 872 AN22JI3VX1 $T=297920 33600 0 0 $X=297490 $Y=32960
X9540 1364 1362 1116 1115 880 547 897 AN22JI3VX1 $T=344960 168000 1 180 $X=340610 $Y=167360
X9541 1364 1362 604 609 920 613 619 AN22JI3VX1 $T=380240 132160 0 0 $X=379810 $Y=131520
X9542 1364 1362 604 612 625 624 619 AN22JI3VX1 $T=383040 141120 1 0 $X=382610 $Y=136000
X9543 1364 1362 623 920 620 615 618 AN22JI3VX1 $T=389760 123200 1 180 $X=385410 $Y=122560
X9544 1364 1362 480 486 659 NO2JI3VX2 $T=301280 123200 1 180 $X=296370 $Y=122560
X9545 1364 1362 140 132 1178 967 AO21JI3VX1 $T=80640 194880 1 0 $X=80210 $Y=189760
X9546 1364 1362 776 761 1002 1193 AO21JI3VX1 $T=146720 123200 0 180 $X=141810 $Y=118080
X9547 1364 1362 1431 1022 323 1388 AO21JI3VX1 $T=186480 176960 0 0 $X=186050 $Y=176320
X9548 1364 1362 377 1239 53 373 AO21JI3VX1 $T=240240 194880 1 180 $X=235330 $Y=194240
X9549 1364 1362 545 530 877 542 AO21JI3VX1 $T=327040 185920 1 0 $X=326610 $Y=180800
X9550 1364 1362 567 892 1158 1116 AO21JI3VX1 $T=348320 159040 1 180 $X=343410 $Y=158400
X9551 1364 1362 902 530 877 588 AO21JI3VX1 $T=345520 185920 1 0 $X=345090 $Y=180800
X9552 1364 1362 384 616 553 918 AO21JI3VX1 $T=375760 159040 1 0 $X=375330 $Y=153920
X9553 1364 1362 486 32 480 NA2I1JI3VX2 $T=300720 105280 0 0 $X=300290 $Y=104640
X9554 1364 1362 480 30 1104 NA2I1JI3VX2 $T=313040 123200 0 0 $X=312610 $Y=122560
X9555 1364 1362 946 70 enable 87 NA22JI3VX1 $T=40880 176960 1 0 $X=40450 $Y=171840
X9556 1364 1362 111 706 92 707 NA22JI3VX1 $T=61040 176960 0 180 $X=56690 $Y=171840
X9557 1364 1362 290 240 315 1415 NA22JI3VX1 $T=179200 176960 1 0 $X=178770 $Y=171840
X9558 1364 1362 349 246 664 1050 NA22JI3VX1 $T=204400 203840 1 0 $X=203970 $Y=198720
X9559 1364 1362 414 1082 411 408 NA22JI3VX1 $T=258720 176960 1 180 $X=254370 $Y=176320
X9560 1364 1362 855 1153 858 449 NA22JI3VX1 $T=271040 185920 0 0 $X=270610 $Y=185280
X9561 1364 1362 1119 21 897 58 NA22JI3VX1 $T=348880 168000 0 0 $X=348450 $Y=167360
X9562 1364 1362 620 636 1147 25 NA22JI3VX1 $T=394800 105280 0 0 $X=394370 $Y=104640
X9563 1364 1362 384 1244 409 531 MU2JI3VX0 $T=250320 24640 0 0 $X=249890 $Y=24000
X9564 1364 1362 384 608 592 643 MU2JI3VX0 $T=380240 24640 0 0 $X=379810 $Y=24000
X9565 1364 1362 384 927 640 597 MU2JI3VX0 $T=402640 24640 1 180 $X=396610 $Y=24000
X9566 1364 1362 384 932 930 1140 MU2JI3VX0 $T=408240 33600 0 180 $X=402210 $Y=28480
X9567 1364 1362 306 365 141 313 OR3JI3VX1 $T=188160 33600 1 0 $X=187730 $Y=28480
X9568 1364 1362 334 1334 799 808 OR3JI3VX1 $T=202720 194880 1 0 $X=202290 $Y=189760
X9569 1364 1362 438 416 1080 851 OR3JI3VX1 $T=258720 168000 0 0 $X=258290 $Y=167360
X9570 1364 1362 851 1393 849 1432 OR3JI3VX1 $T=263200 168000 0 180 $X=258850 $Y=162880
X9571 1364 1362 876 577 887 1117 OR3JI3VX1 $T=350000 33600 0 180 $X=345650 $Y=28480
X9572 1364 1362 131 704 94 1163 702 ON211JI3VX1 $T=49840 159040 1 0 $X=49410 $Y=153920
X9573 1364 1362 90 2 1300 1302 705 ON211JI3VX1 $T=54320 168000 0 0 $X=53890 $Y=167360
X9574 1364 1362 133 1397 134 1174 959 ON211JI3VX1 $T=72800 176960 0 180 $X=68450 $Y=171840
X9575 1364 1362 242 1006 281 1001 1007 ON211JI3VX1 $T=154000 114240 1 0 $X=153570 $Y=109120
X9576 1364 1362 281 782 784 1308 273 ON211JI3VX1 $T=166880 114240 0 0 $X=166450 $Y=113600
X9577 1364 1362 281 794 783 1213 1025 ON211JI3VX1 $T=178080 123200 1 0 $X=177650 $Y=118080
X9578 1364 1362 798 799 300 11 800 ON211JI3VX1 $T=190960 194880 0 0 $X=190530 $Y=194240
X9579 1364 1362 308 801 310 1032 803 ON211JI3VX1 $T=191520 203840 1 0 $X=191090 $Y=198720
X9580 1364 1362 1226 48 800 801 1037 ON211JI3VX1 $T=196000 194880 0 0 $X=195570 $Y=194240
X9581 1364 1362 323 317 42 356 332 ON211JI3VX1 $T=198800 176960 0 0 $X=198370 $Y=176320
X9582 1364 1362 347 1357 806 1229 1230 ON211JI3VX1 $T=207200 168000 1 0 $X=206770 $Y=162880
X9583 1364 1362 45 1433 355 1053 1434 ON211JI3VX1 $T=218960 159040 0 180 $X=214610 $Y=153920
X9584 1364 1362 140 1234 1336 1053 347 ON211JI3VX1 $T=220640 168000 0 180 $X=216290 $Y=162880
X9585 1364 1362 857 856 1255 1087 435 ON211JI3VX1 $T=273280 176960 0 180 $X=268930 $Y=171840
X9586 1364 1362 619 623 613 1297 607 ON211JI3VX1 $T=385840 132160 1 0 $X=385410 $Y=127040
X9587 1364 1362 1414 70 943 87 AN21JI3VX1 $T=29680 168000 1 0 $X=29250 $Y=162880
X9588 1364 1362 93 949 1300 696 AN21JI3VX1 $T=49840 168000 1 0 $X=49410 $Y=162880
X9589 1364 1362 1165 653 708 707 AN21JI3VX1 $T=56560 176960 0 0 $X=56130 $Y=176320
X9590 1364 1362 118 70 1390 140 AN21JI3VX1 $T=66640 185920 1 180 $X=62850 $Y=185280
X9591 1364 1362 1330 999 239 230 AN21JI3VX1 $T=150080 123200 0 0 $X=149650 $Y=122560
X9592 1364 1362 8 1204 775 247 AN21JI3VX1 $T=154560 123200 0 0 $X=154130 $Y=122560
X9593 1364 1362 791 1215 1411 276 AN21JI3VX1 $T=180880 185920 1 0 $X=180450 $Y=180800
X9594 1364 1362 790 1024 1378 340 AN21JI3VX1 $T=184800 168000 0 0 $X=184370 $Y=167360
X9595 1364 1362 798 1221 1033 333 AN21JI3VX1 $T=194320 194880 0 180 $X=190530 $Y=189760
X9596 1364 1362 1416 1227 43 341 AN21JI3VX1 $T=207200 185920 0 180 $X=203410 $Y=180800
X9597 1364 1362 1045 48 49 13 AN21JI3VX1 $T=210560 194880 0 0 $X=210130 $Y=194240
X9598 1364 1362 1087 820 1336 1044 AN21JI3VX1 $T=216160 168000 0 0 $X=215730 $Y=167360
X9599 1364 1362 1045 1046 1055 1060 AN21JI3VX1 $T=222880 194880 1 180 $X=219090 $Y=194240
X9600 1364 1362 1241 1153 1246 1239 AN21JI3VX1 $T=245840 194880 0 180 $X=242050 $Y=189760
X9601 1364 1362 1069 1071 836 389 AN21JI3VX1 $T=243040 168000 1 0 $X=242610 $Y=162880
X9602 1364 1362 846 410 1075 408 AN21JI3VX1 $T=256480 176960 0 180 $X=252690 $Y=171840
X9603 1364 1362 1251 1083 411 419 AN21JI3VX1 $T=263200 185920 1 180 $X=259410 $Y=185280
X9604 1364 1362 1080 1250 1084 1085 AN21JI3VX1 $T=260400 176960 1 0 $X=259970 $Y=171840
X9605 1364 1362 447 464 1382 456 AN21JI3VX1 $T=281680 185920 0 180 $X=277890 $Y=180800
X9606 1364 1362 1417 1227 877 54 AN21JI3VX1 $T=302960 176960 1 0 $X=302530 $Y=171840
X9607 1364 1362 880 500 54 487 AN21JI3VX1 $T=312480 176960 0 180 $X=308690 $Y=171840
X9608 1364 1362 518 524 1383 543 AN21JI3VX1 $T=322560 168000 1 180 $X=318770 $Y=167360
X9609 1364 1362 523 1107 888 1158 AN21JI3VX1 $T=338240 159040 0 0 $X=337810 $Y=158400
X9610 1364 1362 581 1122 1121 909 AN21JI3VX1 $T=362880 176960 1 180 $X=359090 $Y=176320
X9611 1364 1362 384 616 941 553 AN21JI3VX1 $T=380800 159040 1 0 $X=380370 $Y=153920
X9612 1364 1362 636 620 63 633 AN21JI3VX1 $T=394240 114240 1 0 $X=393810 $Y=109120
X9613 1364 1362 68 945 INJI3VX0 $T=33600 168000 1 0 $X=33170 $Y=162880
X9614 1364 1362 78 69 INJI3VX0 $T=38640 159040 0 180 $X=36530 $Y=153920
X9615 1364 1362 1154 74 INJI3VX0 $T=38640 168000 1 180 $X=36530 $Y=167360
X9616 1364 1362 75 79 INJI3VX0 $T=38640 176960 1 0 $X=38210 $Y=171840
X9617 1364 1362 949 1161 INJI3VX0 $T=47040 168000 1 0 $X=46610 $Y=162880
X9618 1364 1362 700 653 INJI3VX0 $T=52080 185920 0 0 $X=51650 $Y=185280
X9619 1364 1362 96 70 INJI3VX0 $T=56560 176960 1 180 $X=54450 $Y=176320
X9620 1364 1362 113 116 INJI3VX0 $T=63280 150080 1 180 $X=61170 $Y=149440
X9621 1364 1362 122 1171 INJI3VX0 $T=67200 194880 0 180 $X=65090 $Y=189760
X9622 1364 1362 131 1174 INJI3VX0 $T=71680 159040 1 180 $X=69570 $Y=158400
X9623 1364 1362 132 134 INJI3VX0 $T=70560 185920 1 0 $X=70130 $Y=180800
X9624 1364 1362 720 129 INJI3VX0 $T=75040 203840 0 180 $X=72930 $Y=198720
X9625 1364 1362 727 31 INJI3VX0 $T=83440 24640 0 0 $X=83010 $Y=24000
X9626 1364 1362 143 1419 INJI3VX0 $T=84000 33600 0 0 $X=83570 $Y=32960
X9627 1364 1362 709 968 INJI3VX0 $T=94080 24640 1 180 $X=91970 $Y=24000
X9628 1364 1362 733 1418 INJI3VX0 $T=92960 42560 0 0 $X=92530 $Y=41920
X9629 1364 1362 163 736 INJI3VX0 $T=108640 33600 0 180 $X=106530 $Y=28480
X9630 1364 1362 167 743 INJI3VX0 $T=117040 24640 0 0 $X=116610 $Y=24000
X9631 1364 1362 752 977 INJI3VX0 $T=123200 24640 0 0 $X=122770 $Y=24000
X9632 1364 1362 214 760 INJI3VX0 $T=136640 33600 0 0 $X=136210 $Y=32960
X9633 1364 1362 217 761 INJI3VX0 $T=139440 159040 0 0 $X=139010 $Y=158400
X9634 1364 1362 768 1420 INJI3VX0 $T=141680 24640 1 180 $X=139570 $Y=24000
X9635 1364 1362 1002 1330 INJI3VX0 $T=152880 123200 0 180 $X=150770 $Y=118080
X9636 1364 1362 1000 241 INJI3VX0 $T=154560 33600 1 180 $X=152450 $Y=32960
X9637 1364 1362 239 1204 INJI3VX0 $T=152880 123200 1 0 $X=152450 $Y=118080
X9638 1364 1362 298 1368 INJI3VX0 $T=164640 114240 1 180 $X=162530 $Y=113600
X9639 1364 1362 251 1421 INJI3VX0 $T=164640 24640 1 0 $X=164210 $Y=19520
X9640 1364 1362 263 270 INJI3VX0 $T=168000 24640 1 0 $X=167570 $Y=19520
X9641 1364 1362 277 253 INJI3VX0 $T=170800 123200 1 180 $X=168690 $Y=122560
X9642 1364 1362 315 237 INJI3VX0 $T=172480 176960 0 180 $X=170370 $Y=171840
X9643 1364 1362 231 281 INJI3VX0 $T=172480 114240 0 0 $X=172050 $Y=113600
X9644 1364 1362 288 240 INJI3VX0 $T=175840 176960 0 180 $X=173730 $Y=171840
X9645 1364 1362 285 793 INJI3VX0 $T=175840 203840 1 0 $X=175410 $Y=198720
X9646 1364 1362 290 1024 INJI3VX0 $T=178080 168000 0 0 $X=177650 $Y=167360
X9647 1364 1362 1019 300 INJI3VX0 $T=178640 194880 0 0 $X=178210 $Y=194240
X9648 1364 1362 39 1422 INJI3VX0 $T=183120 33600 1 0 $X=182690 $Y=28480
X9649 1364 1362 311 795 INJI3VX0 $T=183680 203840 0 0 $X=183250 $Y=203200
X9650 1364 1362 292 1431 INJI3VX0 $T=184240 176960 0 0 $X=183810 $Y=176320
X9651 1364 1362 798 1387 INJI3VX0 $T=190960 176960 0 0 $X=190530 $Y=176320
X9652 1364 1362 272 1221 INJI3VX0 $T=192080 185920 1 0 $X=191650 $Y=180800
X9653 1364 1362 803 1226 INJI3VX0 $T=204400 203840 0 180 $X=202290 $Y=198720
X9654 1364 1362 43 664 INJI3VX0 $T=203280 194880 0 0 $X=202850 $Y=194240
X9655 1364 1362 346 1042 INJI3VX0 $T=205520 33600 0 0 $X=205090 $Y=32960
X9656 1364 1362 331 345 INJI3VX0 $T=208880 42560 1 180 $X=206770 $Y=41920
X9657 1364 1362 246 1335 INJI3VX0 $T=208320 203840 0 0 $X=207890 $Y=203200
X9658 1364 1362 355 1044 INJI3VX0 $T=209440 176960 1 0 $X=209010 $Y=171840
X9659 1364 1362 349 1046 INJI3VX0 $T=209440 203840 1 0 $X=209010 $Y=198720
X9660 1364 1362 353 1434 INJI3VX0 $T=211120 159040 1 0 $X=210690 $Y=153920
X9661 1364 1362 492 1053 INJI3VX0 $T=215040 168000 1 0 $X=214610 $Y=162880
X9662 1364 1362 1045 50 INJI3VX0 $T=215600 185920 0 0 $X=215170 $Y=185280
X9663 1364 1362 390 807 INJI3VX0 $T=219520 185920 1 180 $X=217410 $Y=185280
X9664 1364 1362 364 1423 INJI3VX0 $T=219520 33600 1 0 $X=219090 $Y=28480
X9665 1364 1362 399 1316 INJI3VX0 $T=233520 33600 0 180 $X=231410 $Y=28480
X9666 1364 1362 1065 834 INJI3VX0 $T=241920 185920 0 0 $X=241490 $Y=185280
X9667 1364 1362 409 1424 INJI3VX0 $T=246960 24640 1 180 $X=244850 $Y=24000
X9668 1364 1362 839 385 INJI3VX0 $T=250320 185920 0 180 $X=248210 $Y=180800
X9669 1364 1362 393 410 INJI3VX0 $T=257040 185920 1 180 $X=254930 $Y=185280
X9670 1364 1362 408 1250 INJI3VX0 $T=257600 176960 1 0 $X=257170 $Y=171840
X9671 1364 1362 417 1082 INJI3VX0 $T=262640 194880 0 180 $X=260530 $Y=189760
X9672 1364 1362 423 1153 INJI3VX0 $T=264320 194880 0 180 $X=262210 $Y=189760
X9673 1364 1362 854 419 INJI3VX0 $T=265440 185920 0 180 $X=263330 $Y=180800
X9674 1364 1362 428 1083 INJI3VX0 $T=266000 194880 0 180 $X=263890 $Y=189760
X9675 1364 1362 17 431 INJI3VX0 $T=267680 194880 0 180 $X=265570 $Y=189760
X9676 1364 1362 437 1425 INJI3VX0 $T=269360 24640 1 180 $X=267250 $Y=24000
X9677 1364 1362 858 1239 INJI3VX0 $T=273280 194880 0 180 $X=271170 $Y=189760
X9678 1364 1362 441 1089 INJI3VX0 $T=272160 42560 0 0 $X=271730 $Y=41920
X9679 1364 1362 453 1426 INJI3VX0 $T=276640 33600 0 0 $X=276210 $Y=32960
X9680 1364 1362 855 464 INJI3VX0 $T=278880 185920 0 0 $X=278450 $Y=185280
X9681 1364 1362 872 1099 INJI3VX0 $T=295120 42560 0 0 $X=294690 $Y=41920
X9682 1364 1362 482 873 INJI3VX0 $T=297360 168000 1 0 $X=296930 $Y=162880
X9683 1364 1362 475 1427 INJI3VX0 $T=300720 24640 0 180 $X=298610 $Y=19520
X9684 1364 1362 55 510 INJI3VX0 $T=315280 33600 0 0 $X=314850 $Y=32960
X9685 1364 1362 1096 1107 INJI3VX0 $T=319760 159040 0 0 $X=319330 $Y=158400
X9686 1364 1362 532 884 INJI3VX0 $T=321440 168000 0 180 $X=319330 $Y=162880
X9687 1364 1362 1109 1108 INJI3VX0 $T=323680 24640 1 180 $X=321570 $Y=24000
X9688 1364 1362 537 890 INJI3VX0 $T=333760 33600 1 0 $X=333330 $Y=28480
X9689 1364 1362 57 556 INJI3VX0 $T=337680 176960 0 0 $X=337250 $Y=176320
X9690 1364 1362 58 1115 INJI3VX0 $T=340480 176960 1 0 $X=340050 $Y=171840
X9691 1364 1362 1122 902 INJI3VX0 $T=344400 185920 0 0 $X=343970 $Y=185280
X9692 1364 1362 530 903 INJI3VX0 $T=345520 194880 1 0 $X=345090 $Y=189760
X9693 1364 1362 567 562 INJI3VX0 $T=347760 168000 0 180 $X=345650 $Y=162880
X9694 1364 1362 1128 568 INJI3VX0 $T=346640 51520 1 0 $X=346210 $Y=46400
X9695 1364 1362 575 571 INJI3VX0 $T=347760 176960 1 0 $X=347330 $Y=171840
X9696 1364 1362 566 563 INJI3VX0 $T=348320 212800 1 0 $X=347890 $Y=207680
X9697 1364 1362 581 21 INJI3VX0 $T=362880 176960 0 180 $X=360770 $Y=171840
X9698 1364 1362 909 1123 INJI3VX0 $T=364560 176960 1 180 $X=362450 $Y=176320
X9699 1364 1362 61 1428 INJI3VX0 $T=367920 33600 1 180 $X=365810 $Y=32960
X9700 1364 1362 592 593 INJI3VX0 $T=374640 24640 0 0 $X=374210 $Y=24000
X9701 1364 1362 595 1294 INJI3VX0 $T=375200 42560 1 0 $X=374770 $Y=37440
X9702 1364 1362 606 612 INJI3VX0 $T=381360 141120 0 180 $X=379250 $Y=136000
X9703 1364 1362 615 609 INJI3VX0 $T=384160 123200 1 180 $X=382050 $Y=122560
X9704 1364 1362 604 618 INJI3VX0 $T=385840 132160 0 0 $X=385410 $Y=131520
X9705 1364 1362 639 1297 INJI3VX0 $T=389200 123200 1 0 $X=388770 $Y=118080
X9706 1364 1362 1139 624 INJI3VX0 $T=390880 150080 1 180 $X=388770 $Y=149440
X9707 1364 1362 633 1147 INJI3VX0 $T=392560 123200 0 0 $X=392130 $Y=122560
X9708 1364 1362 1146 631 INJI3VX0 $T=394240 159040 1 180 $X=392130 $Y=158400
X9709 1364 1362 640 1429 INJI3VX0 $T=397040 24640 1 180 $X=394930 $Y=24000
X9710 1364 1362 628 925 INJI3VX0 $T=395920 159040 1 0 $X=395490 $Y=153920
X9711 1364 1362 1413 634 INJI3VX0 $T=398160 141120 0 180 $X=396050 $Y=136000
X9712 1364 1362 930 630 INJI3VX0 $T=405440 33600 1 180 $X=403330 $Y=32960
X9713 1364 1362 708 1370 696 114 NO3I1JI3VX1 $T=57120 168000 1 0 $X=56690 $Y=162880
X9714 1364 1362 791 1412 40 1031 NO3I1JI3VX1 $T=187040 185920 1 0 $X=186610 $Y=180800
X9715 1364 1362 1229 212 231 1433 NO3I1JI3VX1 $T=206080 159040 0 180 $X=201170 $Y=153920
X9716 1364 1362 1075 820 407 1432 NO3I1JI3VX1 $T=254240 168000 1 0 $X=253810 $Y=162880
X9717 1364 1362 518 1396 881 507 NO3I1JI3VX1 $T=319760 168000 0 180 $X=314850 $Y=162880
X9718 1364 1362 DECAP25JI3V $T=20160 24640 1 0 $X=19730 $Y=19520
X9719 1364 1362 DECAP25JI3V $T=20160 24640 0 0 $X=19730 $Y=24000
X9720 1364 1362 DECAP25JI3V $T=20160 33600 1 0 $X=19730 $Y=28480
X9721 1364 1362 DECAP25JI3V $T=20160 42560 1 0 $X=19730 $Y=37440
X9722 1364 1362 DECAP25JI3V $T=20160 42560 0 0 $X=19730 $Y=41920
X9723 1364 1362 DECAP25JI3V $T=20160 51520 1 0 $X=19730 $Y=46400
X9724 1364 1362 DECAP25JI3V $T=20160 51520 0 0 $X=19730 $Y=50880
X9725 1364 1362 DECAP25JI3V $T=20160 60480 1 0 $X=19730 $Y=55360
X9726 1364 1362 DECAP25JI3V $T=20160 60480 0 0 $X=19730 $Y=59840
X9727 1364 1362 DECAP25JI3V $T=20160 69440 1 0 $X=19730 $Y=64320
X9728 1364 1362 DECAP25JI3V $T=20160 69440 0 0 $X=19730 $Y=68800
X9729 1364 1362 DECAP25JI3V $T=20160 78400 1 0 $X=19730 $Y=73280
X9730 1364 1362 DECAP25JI3V $T=20160 78400 0 0 $X=19730 $Y=77760
X9731 1364 1362 DECAP25JI3V $T=20160 87360 1 0 $X=19730 $Y=82240
X9732 1364 1362 DECAP25JI3V $T=20160 87360 0 0 $X=19730 $Y=86720
X9733 1364 1362 DECAP25JI3V $T=20160 96320 1 0 $X=19730 $Y=91200
X9734 1364 1362 DECAP25JI3V $T=20160 141120 0 0 $X=19730 $Y=140480
X9735 1364 1362 DECAP25JI3V $T=20160 194880 0 0 $X=19730 $Y=194240
X9736 1364 1362 DECAP25JI3V $T=20160 203840 1 0 $X=19730 $Y=198720
X9737 1364 1362 DECAP25JI3V $T=20160 203840 0 0 $X=19730 $Y=203200
X9738 1364 1362 DECAP25JI3V $T=20160 212800 1 0 $X=19730 $Y=207680
X9739 1364 1362 DECAP25JI3V $T=20160 212800 0 0 $X=19730 $Y=212160
X9740 1364 1362 DECAP25JI3V $T=34160 33600 1 0 $X=33730 $Y=28480
X9741 1364 1362 DECAP25JI3V $T=34160 60480 0 0 $X=33730 $Y=59840
X9742 1364 1362 DECAP25JI3V $T=34160 87360 0 0 $X=33730 $Y=86720
X9743 1364 1362 DECAP25JI3V $T=34160 203840 1 0 $X=33730 $Y=198720
X9744 1364 1362 DECAP25JI3V $T=34160 212800 1 0 $X=33730 $Y=207680
X9745 1364 1362 DECAP25JI3V $T=34160 212800 0 0 $X=33730 $Y=212160
X9746 1364 1362 DECAP25JI3V $T=48160 87360 0 0 $X=47730 $Y=86720
X9747 1364 1362 DECAP25JI3V $T=48160 212800 0 0 $X=47730 $Y=212160
X9748 1364 1362 DECAP25JI3V $T=57120 132160 0 0 $X=56690 $Y=131520
X9749 1364 1362 DECAP25JI3V $T=80080 123200 1 0 $X=79650 $Y=118080
X9750 1364 1362 DECAP25JI3V $T=85680 96320 0 0 $X=85250 $Y=95680
X9751 1364 1362 DECAP25JI3V $T=86240 87360 0 0 $X=85810 $Y=86720
X9752 1364 1362 DECAP25JI3V $T=86240 105280 1 0 $X=85810 $Y=100160
X9753 1364 1362 DECAP25JI3V $T=89040 114240 0 0 $X=88610 $Y=113600
X9754 1364 1362 DECAP25JI3V $T=93520 105280 0 0 $X=93090 $Y=104640
X9755 1364 1362 DECAP25JI3V $T=110880 87360 0 180 $X=96450 $Y=82240
X9756 1364 1362 DECAP25JI3V $T=215040 114240 0 0 $X=214610 $Y=113600
X9757 1364 1362 DECAP25JI3V $T=223440 123200 0 0 $X=223010 $Y=122560
X9758 1364 1362 DECAP25JI3V $T=231840 96320 1 0 $X=231410 $Y=91200
X9759 1364 1362 DECAP25JI3V $T=257600 114240 0 0 $X=257170 $Y=113600
X9760 1364 1362 DECAP25JI3V $T=271600 114240 0 0 $X=271170 $Y=113600
X9761 1364 1362 DECAP25JI3V $T=295120 78400 0 0 $X=294690 $Y=77760
X9762 1364 1362 DECAP25JI3V $T=308000 132160 0 0 $X=307570 $Y=131520
X9763 1364 1362 DECAP25JI3V $T=312480 105280 0 0 $X=312050 $Y=104640
X9764 1364 1362 DECAP25JI3V $T=313040 194880 0 0 $X=312610 $Y=194240
X9765 1364 1362 DECAP25JI3V $T=318080 123200 0 0 $X=317650 $Y=122560
X9766 1364 1362 DECAP25JI3V $T=333760 114240 1 0 $X=333330 $Y=109120
X9767 1364 1362 DECAP25JI3V $T=336000 105280 1 0 $X=335570 $Y=100160
X9768 1364 1362 DECAP25JI3V $T=338240 87360 1 0 $X=337810 $Y=82240
X9769 1364 1362 DECAP25JI3V $T=350000 212800 1 0 $X=349570 $Y=207680
X9770 1364 1362 DECAP25JI3V $T=351120 203840 0 0 $X=350690 $Y=203200
X9771 1364 1362 DECAP25JI3V $T=352240 212800 0 0 $X=351810 $Y=212160
X9772 1364 1362 DECAP25JI3V $T=352800 203840 1 0 $X=352370 $Y=198720
X9773 1364 1362 DECAP25JI3V $T=364000 212800 1 0 $X=363570 $Y=207680
X9774 1364 1362 DECAP25JI3V $T=365120 203840 0 0 $X=364690 $Y=203200
X9775 1364 1362 DECAP25JI3V $T=366240 212800 0 0 $X=365810 $Y=212160
X9776 1364 1362 DECAP25JI3V $T=366800 203840 1 0 $X=366370 $Y=198720
X9777 1364 1362 DECAP25JI3V $T=370160 194880 1 0 $X=369730 $Y=189760
X9778 1364 1362 DECAP25JI3V $T=371280 194880 0 0 $X=370850 $Y=194240
X9779 1364 1362 DECAP25JI3V $T=378000 212800 1 0 $X=377570 $Y=207680
X9780 1364 1362 DECAP25JI3V $T=379120 185920 0 0 $X=378690 $Y=185280
X9781 1364 1362 DECAP25JI3V $T=379120 203840 0 0 $X=378690 $Y=203200
X9782 1364 1362 DECAP25JI3V $T=380240 212800 0 0 $X=379810 $Y=212160
X9783 1364 1362 DECAP25JI3V $T=380800 176960 0 0 $X=380370 $Y=176320
X9784 1364 1362 DECAP25JI3V $T=380800 203840 1 0 $X=380370 $Y=198720
X9785 1364 1362 DECAP25JI3V $T=381360 176960 1 0 $X=380930 $Y=171840
X9786 1364 1362 DECAP25JI3V $T=384160 194880 1 0 $X=383730 $Y=189760
X9787 1364 1362 DECAP25JI3V $T=385280 194880 0 0 $X=384850 $Y=194240
X9788 1364 1362 DECAP25JI3V $T=389200 185920 1 0 $X=388770 $Y=180800
X9789 1364 1362 DECAP25JI3V $T=392000 212800 1 0 $X=391570 $Y=207680
X9790 1364 1362 DECAP25JI3V $T=393120 185920 0 0 $X=392690 $Y=185280
X9791 1364 1362 DECAP25JI3V $T=393120 203840 0 0 $X=392690 $Y=203200
X9792 1364 1362 DECAP25JI3V $T=394240 212800 0 0 $X=393810 $Y=212160
X9793 1364 1362 DECAP25JI3V $T=394800 176960 0 0 $X=394370 $Y=176320
X9794 1364 1362 DECAP25JI3V $T=394800 203840 1 0 $X=394370 $Y=198720
X9795 1364 1362 DECAP25JI3V $T=395360 176960 1 0 $X=394930 $Y=171840
X9796 1364 1362 DECAP25JI3V $T=398160 194880 1 0 $X=397730 $Y=189760
X9797 1364 1362 DECAP25JI3V $T=398720 141120 0 0 $X=398290 $Y=140480
X9798 1364 1362 DECAP25JI3V $T=398720 150080 1 0 $X=398290 $Y=144960
X9799 1364 1362 DECAP25JI3V $T=399280 194880 0 0 $X=398850 $Y=194240
X9800 1364 1362 DECAP25JI3V $T=399840 159040 0 0 $X=399410 $Y=158400
X9801 1364 1362 DECAP25JI3V $T=400400 78400 0 0 $X=399970 $Y=77760
X9802 1364 1362 DECAP25JI3V $T=400400 96320 0 0 $X=399970 $Y=95680
X9803 1364 1362 DECAP25JI3V $T=414400 168000 0 180 $X=399970 $Y=162880
X9804 1364 1362 DECAP25JI3V $T=402080 141120 1 0 $X=401650 $Y=136000
X9805 1364 1362 DECAP25JI3V $T=403200 185920 1 0 $X=402770 $Y=180800
X9806 1364 1362 DECAP25JI3V $T=404320 159040 1 0 $X=403890 $Y=153920
X9807 1364 1362 DECAP25JI3V $T=406000 24640 1 0 $X=405570 $Y=19520
X9808 1364 1362 DECAP25JI3V $T=406000 212800 1 0 $X=405570 $Y=207680
X9809 1364 1362 DECAP25JI3V $T=406560 105280 0 0 $X=406130 $Y=104640
X9810 1364 1362 DECAP25JI3V $T=406560 114240 1 0 $X=406130 $Y=109120
X9811 1364 1362 DECAP25JI3V $T=407120 185920 0 0 $X=406690 $Y=185280
X9812 1364 1362 DECAP25JI3V $T=407120 203840 0 0 $X=406690 $Y=203200
X9813 1364 1362 DECAP25JI3V $T=407680 168000 0 0 $X=407250 $Y=167360
X9814 1364 1362 DECAP25JI3V $T=408800 150080 0 0 $X=408370 $Y=149440
X9815 1364 1362 DECAP25JI3V $T=408800 176960 0 0 $X=408370 $Y=176320
X9816 1364 1362 DECAP25JI3V $T=408800 203840 1 0 $X=408370 $Y=198720
X9817 1364 1362 DECAP25JI3V $T=409360 24640 0 0 $X=408930 $Y=24000
X9818 1364 1362 DECAP25JI3V $T=409360 176960 1 0 $X=408930 $Y=171840
X9819 1364 1362 DECAP25JI3V $T=409920 132160 1 0 $X=409490 $Y=127040
X9820 1364 1362 DECAP25JI3V $T=412720 132160 0 0 $X=412290 $Y=131520
X9821 1364 1362 DECAP25JI3V $T=412720 141120 0 0 $X=412290 $Y=140480
X9822 1364 1362 DECAP25JI3V $T=412720 150080 1 0 $X=412290 $Y=144960
X9823 1364 1362 DECAP25JI3V $T=413280 42560 1 0 $X=412850 $Y=37440
X9824 1364 1362 DECAP25JI3V $T=413280 60480 0 0 $X=412850 $Y=59840
X9825 1364 1362 DECAP25JI3V $T=413280 69440 1 0 $X=412850 $Y=64320
X9826 1364 1362 DECAP25JI3V $T=413280 69440 0 0 $X=412850 $Y=68800
X9827 1364 1362 DECAP25JI3V $T=413280 105280 1 0 $X=412850 $Y=100160
X9828 1364 1362 DECAP25JI3V $T=413280 194880 0 0 $X=412850 $Y=194240
X9829 1364 1362 DECAP25JI3V $T=414400 78400 0 0 $X=413970 $Y=77760
X9830 1364 1362 DECAP25JI3V $T=414400 96320 0 0 $X=413970 $Y=95680
X9831 1364 1362 DECAP25JI3V $T=414400 168000 1 0 $X=413970 $Y=162880
X9832 1364 1362 DECAP25JI3V $T=417200 185920 1 0 $X=416770 $Y=180800
X9833 1364 1362 DECAP25JI3V $T=418320 159040 1 0 $X=417890 $Y=153920
X9834 1364 1362 DECAP25JI3V $T=421120 185920 0 0 $X=420690 $Y=185280
X9835 1364 1362 DECAP25JI3V $T=421120 203840 0 0 $X=420690 $Y=203200
X9836 1364 1362 DECAP15JI3V $T=20160 33600 0 0 $X=19730 $Y=32960
X9837 1364 1362 DECAP15JI3V $T=20160 96320 0 0 $X=19730 $Y=95680
X9838 1364 1362 DECAP15JI3V $T=20160 141120 1 0 $X=19730 $Y=136000
X9839 1364 1362 DECAP15JI3V $T=34160 24640 1 0 $X=33730 $Y=19520
X9840 1364 1362 DECAP15JI3V $T=34160 60480 1 0 $X=33730 $Y=55360
X9841 1364 1362 DECAP15JI3V $T=34160 69440 0 0 $X=33730 $Y=68800
X9842 1364 1362 DECAP15JI3V $T=34160 78400 1 0 $X=33730 $Y=73280
X9843 1364 1362 DECAP15JI3V $T=34160 203840 0 0 $X=33730 $Y=203200
X9844 1364 1362 DECAP15JI3V $T=48160 60480 0 0 $X=47730 $Y=59840
X9845 1364 1362 DECAP15JI3V $T=48160 212800 1 0 $X=47730 $Y=207680
X9846 1364 1362 DECAP15JI3V $T=54880 114240 0 0 $X=54450 $Y=113600
X9847 1364 1362 DECAP15JI3V $T=61040 69440 1 0 $X=60610 $Y=64320
X9848 1364 1362 DECAP15JI3V $T=62720 69440 0 0 $X=62290 $Y=68800
X9849 1364 1362 DECAP15JI3V $T=62720 78400 1 0 $X=62290 $Y=73280
X9850 1364 1362 DECAP15JI3V $T=80080 132160 1 0 $X=79650 $Y=127040
X9851 1364 1362 DECAP15JI3V $T=84000 123200 0 0 $X=83570 $Y=122560
X9852 1364 1362 DECAP15JI3V $T=86800 96320 1 0 $X=86370 $Y=91200
X9853 1364 1362 DECAP15JI3V $T=90160 185920 1 0 $X=89730 $Y=180800
X9854 1364 1362 DECAP15JI3V $T=90160 212800 1 0 $X=89730 $Y=207680
X9855 1364 1362 DECAP15JI3V $T=91280 150080 0 0 $X=90850 $Y=149440
X9856 1364 1362 DECAP15JI3V $T=91840 159040 1 0 $X=91410 $Y=153920
X9857 1364 1362 DECAP15JI3V $T=94080 123200 1 0 $X=93650 $Y=118080
X9858 1364 1362 DECAP15JI3V $T=95200 69440 0 0 $X=94770 $Y=68800
X9859 1364 1362 DECAP15JI3V $T=99680 96320 0 0 $X=99250 $Y=95680
X9860 1364 1362 DECAP15JI3V $T=100240 78400 0 0 $X=99810 $Y=77760
X9861 1364 1362 DECAP15JI3V $T=103040 114240 0 0 $X=102610 $Y=113600
X9862 1364 1362 DECAP15JI3V $T=108080 96320 0 0 $X=107650 $Y=95680
X9863 1364 1362 DECAP15JI3V $T=123200 78400 1 0 $X=122770 $Y=73280
X9864 1364 1362 DECAP15JI3V $T=128240 194880 1 0 $X=127810 $Y=189760
X9865 1364 1362 DECAP15JI3V $T=137760 159040 1 180 $X=128930 $Y=158400
X9866 1364 1362 DECAP15JI3V $T=131600 78400 0 0 $X=131170 $Y=77760
X9867 1364 1362 DECAP15JI3V $T=151200 168000 1 0 $X=150770 $Y=162880
X9868 1364 1362 DECAP15JI3V $T=162960 78400 0 0 $X=162530 $Y=77760
X9869 1364 1362 DECAP15JI3V $T=210000 87360 1 0 $X=209570 $Y=82240
X9870 1364 1362 DECAP15JI3V $T=215600 42560 0 0 $X=215170 $Y=41920
X9871 1364 1362 DECAP15JI3V $T=215600 51520 1 0 $X=215170 $Y=46400
X9872 1364 1362 DECAP15JI3V $T=223440 33600 0 0 $X=223010 $Y=32960
X9873 1364 1362 DECAP15JI3V $T=223440 69440 0 0 $X=223010 $Y=68800
X9874 1364 1362 DECAP15JI3V $T=223440 78400 1 0 $X=223010 $Y=73280
X9875 1364 1362 DECAP15JI3V $T=223440 96320 1 0 $X=223010 $Y=91200
X9876 1364 1362 DECAP15JI3V $T=223440 105280 1 0 $X=223010 $Y=100160
X9877 1364 1362 DECAP15JI3V $T=223440 114240 1 0 $X=223010 $Y=109120
X9878 1364 1362 DECAP15JI3V $T=229040 114240 0 0 $X=228610 $Y=113600
X9879 1364 1362 DECAP15JI3V $T=258720 78400 0 0 $X=258290 $Y=77760
X9880 1364 1362 DECAP15JI3V $T=267120 212800 1 0 $X=266690 $Y=207680
X9881 1364 1362 DECAP15JI3V $T=268800 212800 0 0 $X=268370 $Y=212160
X9882 1364 1362 DECAP15JI3V $T=276640 105280 1 0 $X=276210 $Y=100160
X9883 1364 1362 DECAP15JI3V $T=279440 42560 0 0 $X=279010 $Y=41920
X9884 1364 1362 DECAP15JI3V $T=280560 185920 0 0 $X=280130 $Y=185280
X9885 1364 1362 DECAP15JI3V $T=294560 96320 0 0 $X=294130 $Y=95680
X9886 1364 1362 DECAP15JI3V $T=298480 194880 1 0 $X=298050 $Y=189760
X9887 1364 1362 DECAP15JI3V $T=300720 114240 1 0 $X=300290 $Y=109120
X9888 1364 1362 DECAP15JI3V $T=327600 203840 0 0 $X=327170 $Y=203200
X9889 1364 1362 DECAP15JI3V $T=336000 96320 0 0 $X=335570 $Y=95680
X9890 1364 1362 DECAP15JI3V $T=337120 96320 1 0 $X=336690 $Y=91200
X9891 1364 1362 DECAP15JI3V $T=337120 114240 0 0 $X=336690 $Y=113600
X9892 1364 1362 DECAP15JI3V $T=344960 194880 0 0 $X=344530 $Y=194240
X9893 1364 1362 DECAP15JI3V $T=350000 105280 1 0 $X=349570 $Y=100160
X9894 1364 1362 DECAP15JI3V $T=350000 185920 1 0 $X=349570 $Y=180800
X9895 1364 1362 DECAP15JI3V $T=351680 51520 1 0 $X=351250 $Y=46400
X9896 1364 1362 DECAP15JI3V $T=351680 69440 0 0 $X=351250 $Y=68800
X9897 1364 1362 DECAP15JI3V $T=351680 78400 1 0 $X=351250 $Y=73280
X9898 1364 1362 DECAP15JI3V $T=352240 24640 0 0 $X=351810 $Y=24000
X9899 1364 1362 DECAP15JI3V $T=381920 141120 1 180 $X=373090 $Y=140480
X9900 1364 1362 DECAP15JI3V $T=388640 96320 0 180 $X=379810 $Y=91200
X9901 1364 1362 DECAP15JI3V $T=380800 185920 1 0 $X=380370 $Y=180800
X9902 1364 1362 DECAP15JI3V $T=381360 78400 1 0 $X=380930 $Y=73280
X9903 1364 1362 DECAP15JI3V $T=416640 33600 0 180 $X=407810 $Y=28480
X9904 1364 1362 DECAP15JI3V $T=408240 212800 0 0 $X=407810 $Y=212160
X9905 1364 1362 DECAP15JI3V $T=411040 114240 0 0 $X=410610 $Y=113600
X9906 1364 1362 DECAP15JI3V $T=412160 194880 1 0 $X=411730 $Y=189760
X9907 1364 1362 DECAP15JI3V $T=413280 33600 0 0 $X=412850 $Y=32960
X9908 1364 1362 DECAP15JI3V $T=413280 60480 1 0 $X=412850 $Y=55360
X9909 1364 1362 DECAP15JI3V $T=416080 123200 1 0 $X=415650 $Y=118080
X9910 1364 1362 DECAP15JI3V $T=416080 141120 1 0 $X=415650 $Y=136000
X9911 1364 1362 DECAP15JI3V $T=418880 42560 0 0 $X=418450 $Y=41920
X9912 1364 1362 DECAP15JI3V $T=418880 51520 1 0 $X=418450 $Y=46400
X9913 1364 1362 DECAP15JI3V $T=418880 51520 0 0 $X=418450 $Y=50880
X9914 1364 1362 DECAP15JI3V $T=420000 24640 1 0 $X=419570 $Y=19520
X9915 1364 1362 DECAP15JI3V $T=420000 212800 1 0 $X=419570 $Y=207680
X9916 1364 1362 DECAP15JI3V $T=422800 150080 0 0 $X=422370 $Y=149440
X9917 1364 1362 DECAP15JI3V $T=422800 176960 0 0 $X=422370 $Y=176320
X9918 1364 1362 DECAP15JI3V $T=422800 203840 1 0 $X=422370 $Y=198720
X9919 1364 1362 DECAP15JI3V $T=423920 132160 1 0 $X=423490 $Y=127040
X9920 1364 1362 DECAP15JI3V $T=426720 132160 0 0 $X=426290 $Y=131520
X9921 1364 1362 DECAP15JI3V $T=426720 141120 0 0 $X=426290 $Y=140480
X9922 1364 1362 DECAP15JI3V $T=426720 150080 1 0 $X=426290 $Y=144960
X9923 1364 1362 DECAP7JI3V $T=20160 105280 1 0 $X=19730 $Y=100160
X9924 1364 1362 DECAP7JI3V $T=20160 150080 0 0 $X=19730 $Y=149440
X9925 1364 1362 DECAP7JI3V $T=20160 168000 1 0 $X=19730 $Y=162880
X9926 1364 1362 DECAP7JI3V $T=20160 168000 0 0 $X=19730 $Y=167360
X9927 1364 1362 DECAP7JI3V $T=25760 114240 0 0 $X=25330 $Y=113600
X9928 1364 1362 DECAP7JI3V $T=25760 123200 1 0 $X=25330 $Y=118080
X9929 1364 1362 DECAP7JI3V $T=25760 176960 0 0 $X=25330 $Y=176320
X9930 1364 1362 DECAP7JI3V $T=28560 33600 0 0 $X=28130 $Y=32960
X9931 1364 1362 DECAP7JI3V $T=28560 96320 0 0 $X=28130 $Y=95680
X9932 1364 1362 DECAP7JI3V $T=32480 33600 0 0 $X=32050 $Y=32960
X9933 1364 1362 DECAP7JI3V $T=34160 42560 1 0 $X=33730 $Y=37440
X9934 1364 1362 DECAP7JI3V $T=34160 42560 0 0 $X=33730 $Y=41920
X9935 1364 1362 DECAP7JI3V $T=34160 51520 1 0 $X=33730 $Y=46400
X9936 1364 1362 DECAP7JI3V $T=34160 51520 0 0 $X=33730 $Y=50880
X9937 1364 1362 DECAP7JI3V $T=34160 69440 1 0 $X=33730 $Y=64320
X9938 1364 1362 DECAP7JI3V $T=34160 78400 0 0 $X=33730 $Y=77760
X9939 1364 1362 DECAP7JI3V $T=34160 96320 1 0 $X=33730 $Y=91200
X9940 1364 1362 DECAP7JI3V $T=36400 33600 0 0 $X=35970 $Y=32960
X9941 1364 1362 DECAP7JI3V $T=36960 123200 1 0 $X=36530 $Y=118080
X9942 1364 1362 DECAP7JI3V $T=38080 42560 1 0 $X=37650 $Y=37440
X9943 1364 1362 DECAP7JI3V $T=38080 42560 0 0 $X=37650 $Y=41920
X9944 1364 1362 DECAP7JI3V $T=38080 51520 1 0 $X=37650 $Y=46400
X9945 1364 1362 DECAP7JI3V $T=38080 51520 0 0 $X=37650 $Y=50880
X9946 1364 1362 DECAP7JI3V $T=38080 69440 1 0 $X=37650 $Y=64320
X9947 1364 1362 DECAP7JI3V $T=38080 96320 1 0 $X=37650 $Y=91200
X9948 1364 1362 DECAP7JI3V $T=39760 24640 0 0 $X=39330 $Y=24000
X9949 1364 1362 DECAP7JI3V $T=39760 194880 0 0 $X=39330 $Y=194240
X9950 1364 1362 DECAP7JI3V $T=40320 33600 0 0 $X=39890 $Y=32960
X9951 1364 1362 DECAP7JI3V $T=42000 69440 1 0 $X=41570 $Y=64320
X9952 1364 1362 DECAP7JI3V $T=42560 24640 1 0 $X=42130 $Y=19520
X9953 1364 1362 DECAP7JI3V $T=42560 203840 0 0 $X=42130 $Y=203200
X9954 1364 1362 DECAP7JI3V $T=43680 24640 0 0 $X=43250 $Y=24000
X9955 1364 1362 DECAP7JI3V $T=43680 194880 0 0 $X=43250 $Y=194240
X9956 1364 1362 DECAP7JI3V $T=46480 24640 1 0 $X=46050 $Y=19520
X9957 1364 1362 DECAP7JI3V $T=46480 203840 0 0 $X=46050 $Y=203200
X9958 1364 1362 DECAP7JI3V $T=47600 24640 0 0 $X=47170 $Y=24000
X9959 1364 1362 DECAP7JI3V $T=50400 24640 1 0 $X=49970 $Y=19520
X9960 1364 1362 DECAP7JI3V $T=50400 203840 0 0 $X=49970 $Y=203200
X9961 1364 1362 DECAP7JI3V $T=51520 24640 0 0 $X=51090 $Y=24000
X9962 1364 1362 DECAP7JI3V $T=54320 203840 0 0 $X=53890 $Y=203200
X9963 1364 1362 DECAP7JI3V $T=56560 60480 0 0 $X=56130 $Y=59840
X9964 1364 1362 DECAP7JI3V $T=56560 212800 1 0 $X=56130 $Y=207680
X9965 1364 1362 DECAP7JI3V $T=59920 51520 0 0 $X=59490 $Y=50880
X9966 1364 1362 DECAP7JI3V $T=60480 212800 1 0 $X=60050 $Y=207680
X9967 1364 1362 DECAP7JI3V $T=62160 212800 0 0 $X=61730 $Y=212160
X9968 1364 1362 DECAP7JI3V $T=62720 194880 0 0 $X=62290 $Y=194240
X9969 1364 1362 DECAP7JI3V $T=63280 114240 1 0 $X=62850 $Y=109120
X9970 1364 1362 DECAP7JI3V $T=64400 212800 1 0 $X=63970 $Y=207680
X9971 1364 1362 DECAP7JI3V $T=66080 212800 0 0 $X=65650 $Y=212160
X9972 1364 1362 DECAP7JI3V $T=67200 114240 1 0 $X=66770 $Y=109120
X9973 1364 1362 DECAP7JI3V $T=68320 212800 1 0 $X=67890 $Y=207680
X9974 1364 1362 DECAP7JI3V $T=70000 212800 0 0 $X=69570 $Y=212160
X9975 1364 1362 DECAP7JI3V $T=71120 78400 1 0 $X=70690 $Y=73280
X9976 1364 1362 DECAP7JI3V $T=71120 114240 1 0 $X=70690 $Y=109120
X9977 1364 1362 DECAP7JI3V $T=71120 132160 0 0 $X=70690 $Y=131520
X9978 1364 1362 DECAP7JI3V $T=80640 185920 0 0 $X=80210 $Y=185280
X9979 1364 1362 DECAP7JI3V $T=88480 132160 1 0 $X=88050 $Y=127040
X9980 1364 1362 DECAP7JI3V $T=90720 194880 0 0 $X=90290 $Y=194240
X9981 1364 1362 DECAP7JI3V $T=91280 185920 0 0 $X=90850 $Y=185280
X9982 1364 1362 DECAP7JI3V $T=92400 123200 0 0 $X=91970 $Y=122560
X9983 1364 1362 DECAP7JI3V $T=92400 132160 1 0 $X=91970 $Y=127040
X9984 1364 1362 DECAP7JI3V $T=93520 60480 0 0 $X=93090 $Y=59840
X9985 1364 1362 DECAP7JI3V $T=94640 42560 1 0 $X=94210 $Y=37440
X9986 1364 1362 DECAP7JI3V $T=94640 42560 0 0 $X=94210 $Y=41920
X9987 1364 1362 DECAP7JI3V $T=94640 194880 0 0 $X=94210 $Y=194240
X9988 1364 1362 DECAP7JI3V $T=95200 33600 1 0 $X=94770 $Y=28480
X9989 1364 1362 DECAP7JI3V $T=95200 69440 1 0 $X=94770 $Y=64320
X9990 1364 1362 DECAP7JI3V $T=95200 78400 1 0 $X=94770 $Y=73280
X9991 1364 1362 DECAP7JI3V $T=95200 96320 1 0 $X=94770 $Y=91200
X9992 1364 1362 DECAP7JI3V $T=95200 114240 1 0 $X=94770 $Y=109120
X9993 1364 1362 DECAP7JI3V $T=95200 132160 0 0 $X=94770 $Y=131520
X9994 1364 1362 DECAP7JI3V $T=95200 185920 0 0 $X=94770 $Y=185280
X9995 1364 1362 DECAP7JI3V $T=95200 203840 0 0 $X=94770 $Y=203200
X9996 1364 1362 DECAP7JI3V $T=96320 123200 0 0 $X=95890 $Y=122560
X9997 1364 1362 DECAP7JI3V $T=96320 132160 1 0 $X=95890 $Y=127040
X9998 1364 1362 DECAP7JI3V $T=96320 176960 1 0 $X=95890 $Y=171840
X9999 1364 1362 DECAP7JI3V $T=99120 33600 1 0 $X=98690 $Y=28480
X10000 1364 1362 DECAP7JI3V $T=99120 69440 1 0 $X=98690 $Y=64320
X10001 1364 1362 DECAP7JI3V $T=99120 78400 1 0 $X=98690 $Y=73280
X10002 1364 1362 DECAP7JI3V $T=99120 96320 1 0 $X=98690 $Y=91200
X10003 1364 1362 DECAP7JI3V $T=99120 114240 1 0 $X=98690 $Y=109120
X10004 1364 1362 DECAP7JI3V $T=99120 132160 0 0 $X=98690 $Y=131520
X10005 1364 1362 DECAP7JI3V $T=99120 185920 0 0 $X=98690 $Y=185280
X10006 1364 1362 DECAP7JI3V $T=99120 203840 0 0 $X=98690 $Y=203200
X10007 1364 1362 DECAP7JI3V $T=99680 150080 0 0 $X=99250 $Y=149440
X10008 1364 1362 DECAP7JI3V $T=100240 87360 0 0 $X=99810 $Y=86720
X10009 1364 1362 DECAP7JI3V $T=100240 176960 1 0 $X=99810 $Y=171840
X10010 1364 1362 DECAP7JI3V $T=100800 159040 0 0 $X=100370 $Y=158400
X10011 1364 1362 DECAP7JI3V $T=103040 33600 1 0 $X=102610 $Y=28480
X10012 1364 1362 DECAP7JI3V $T=103040 96320 1 0 $X=102610 $Y=91200
X10013 1364 1362 DECAP7JI3V $T=103040 114240 1 0 $X=102610 $Y=109120
X10014 1364 1362 DECAP7JI3V $T=104160 87360 0 0 $X=103730 $Y=86720
X10015 1364 1362 DECAP7JI3V $T=104720 159040 0 0 $X=104290 $Y=158400
X10016 1364 1362 DECAP7JI3V $T=105840 194880 1 0 $X=105410 $Y=189760
X10017 1364 1362 DECAP7JI3V $T=106960 96320 1 0 $X=106530 $Y=91200
X10018 1364 1362 DECAP7JI3V $T=106960 114240 1 0 $X=106530 $Y=109120
X10019 1364 1362 DECAP7JI3V $T=111440 114240 0 0 $X=111010 $Y=113600
X10020 1364 1362 DECAP7JI3V $T=116480 96320 0 0 $X=116050 $Y=95680
X10021 1364 1362 DECAP7JI3V $T=123200 69440 1 0 $X=122770 $Y=64320
X10022 1364 1362 DECAP7JI3V $T=128240 105280 0 180 $X=123890 $Y=100160
X10023 1364 1362 DECAP7JI3V $T=127120 69440 1 0 $X=126690 $Y=64320
X10024 1364 1362 DECAP7JI3V $T=132160 69440 0 0 $X=131730 $Y=68800
X10025 1364 1362 DECAP7JI3V $T=132160 87360 0 0 $X=131730 $Y=86720
X10026 1364 1362 DECAP7JI3V $T=135520 212800 0 0 $X=135090 $Y=212160
X10027 1364 1362 DECAP7JI3V $T=136080 87360 0 0 $X=135650 $Y=86720
X10028 1364 1362 DECAP7JI3V $T=138320 33600 0 0 $X=137890 $Y=32960
X10029 1364 1362 DECAP7JI3V $T=151760 78400 1 0 $X=151330 $Y=73280
X10030 1364 1362 DECAP7JI3V $T=155680 78400 1 0 $X=155250 $Y=73280
X10031 1364 1362 DECAP7JI3V $T=155680 203840 1 0 $X=155250 $Y=198720
X10032 1364 1362 DECAP7JI3V $T=158480 87360 1 0 $X=158050 $Y=82240
X10033 1364 1362 DECAP7JI3V $T=159600 168000 1 0 $X=159170 $Y=162880
X10034 1364 1362 DECAP7JI3V $T=162400 33600 0 0 $X=161970 $Y=32960
X10035 1364 1362 DECAP7JI3V $T=162960 60480 0 0 $X=162530 $Y=59840
X10036 1364 1362 DECAP7JI3V $T=166320 168000 0 0 $X=165890 $Y=167360
X10037 1364 1362 DECAP7JI3V $T=166880 60480 0 0 $X=166450 $Y=59840
X10038 1364 1362 DECAP7JI3V $T=169680 24640 1 0 $X=169250 $Y=19520
X10039 1364 1362 DECAP7JI3V $T=170240 168000 0 0 $X=169810 $Y=167360
X10040 1364 1362 DECAP7JI3V $T=170800 60480 0 0 $X=170370 $Y=59840
X10041 1364 1362 DECAP7JI3V $T=171360 78400 0 0 $X=170930 $Y=77760
X10042 1364 1362 DECAP7JI3V $T=178080 168000 1 180 $X=173730 $Y=167360
X10043 1364 1362 DECAP7JI3V $T=174720 60480 0 0 $X=174290 $Y=59840
X10044 1364 1362 DECAP7JI3V $T=175280 78400 0 0 $X=174850 $Y=77760
X10045 1364 1362 DECAP7JI3V $T=179200 78400 0 0 $X=178770 $Y=77760
X10046 1364 1362 DECAP7JI3V $T=184240 69440 0 0 $X=183810 $Y=68800
X10047 1364 1362 DECAP7JI3V $T=184800 194880 1 0 $X=184370 $Y=189760
X10048 1364 1362 DECAP7JI3V $T=197680 33600 0 0 $X=197250 $Y=32960
X10049 1364 1362 DECAP7JI3V $T=197680 60480 1 0 $X=197250 $Y=55360
X10050 1364 1362 DECAP7JI3V $T=205520 33600 1 180 $X=201170 $Y=32960
X10051 1364 1362 DECAP7JI3V $T=203280 42560 0 0 $X=202850 $Y=41920
X10052 1364 1362 DECAP7JI3V $T=215040 69440 1 0 $X=214610 $Y=64320
X10053 1364 1362 DECAP7JI3V $T=216160 60480 0 0 $X=215730 $Y=59840
X10054 1364 1362 DECAP7JI3V $T=218400 87360 1 0 $X=217970 $Y=82240
X10055 1364 1362 DECAP7JI3V $T=218960 69440 1 0 $X=218530 $Y=64320
X10056 1364 1362 DECAP7JI3V $T=220080 60480 0 0 $X=219650 $Y=59840
X10057 1364 1362 DECAP7JI3V $T=221200 33600 1 0 $X=220770 $Y=28480
X10058 1364 1362 DECAP7JI3V $T=221200 212800 0 0 $X=220770 $Y=212160
X10059 1364 1362 DECAP7JI3V $T=222320 24640 0 0 $X=221890 $Y=24000
X10060 1364 1362 DECAP7JI3V $T=222320 87360 1 0 $X=221890 $Y=82240
X10061 1364 1362 DECAP7JI3V $T=222880 69440 1 0 $X=222450 $Y=64320
X10062 1364 1362 DECAP7JI3V $T=222880 168000 0 0 $X=222450 $Y=167360
X10063 1364 1362 DECAP7JI3V $T=223440 185920 0 0 $X=223010 $Y=185280
X10064 1364 1362 DECAP7JI3V $T=224000 42560 0 0 $X=223570 $Y=41920
X10065 1364 1362 DECAP7JI3V $T=225120 33600 1 0 $X=224690 $Y=28480
X10066 1364 1362 DECAP7JI3V $T=225120 212800 0 0 $X=224690 $Y=212160
X10067 1364 1362 DECAP7JI3V $T=225680 212800 1 0 $X=225250 $Y=207680
X10068 1364 1362 DECAP7JI3V $T=226240 24640 0 0 $X=225810 $Y=24000
X10069 1364 1362 DECAP7JI3V $T=226240 87360 1 0 $X=225810 $Y=82240
X10070 1364 1362 DECAP7JI3V $T=226800 168000 0 0 $X=226370 $Y=167360
X10071 1364 1362 DECAP7JI3V $T=227360 185920 0 0 $X=226930 $Y=185280
X10072 1364 1362 DECAP7JI3V $T=227920 42560 0 0 $X=227490 $Y=41920
X10073 1364 1362 DECAP7JI3V $T=229040 78400 0 0 $X=228610 $Y=77760
X10074 1364 1362 DECAP7JI3V $T=229040 87360 0 0 $X=228610 $Y=86720
X10075 1364 1362 DECAP7JI3V $T=229040 96320 0 0 $X=228610 $Y=95680
X10076 1364 1362 DECAP7JI3V $T=229040 105280 0 0 $X=228610 $Y=104640
X10077 1364 1362 DECAP7JI3V $T=229040 132160 0 0 $X=228610 $Y=131520
X10078 1364 1362 DECAP7JI3V $T=231840 78400 1 0 $X=231410 $Y=73280
X10079 1364 1362 DECAP7JI3V $T=231840 123200 1 0 $X=231410 $Y=118080
X10080 1364 1362 DECAP7JI3V $T=232960 132160 0 0 $X=232530 $Y=131520
X10081 1364 1362 DECAP7JI3V $T=234080 141120 1 0 $X=233650 $Y=136000
X10082 1364 1362 DECAP7JI3V $T=235760 78400 1 0 $X=235330 $Y=73280
X10083 1364 1362 DECAP7JI3V $T=235760 123200 1 0 $X=235330 $Y=118080
X10084 1364 1362 DECAP7JI3V $T=239680 78400 1 0 $X=239250 $Y=73280
X10085 1364 1362 DECAP7JI3V $T=243600 78400 1 0 $X=243170 $Y=73280
X10086 1364 1362 DECAP7JI3V $T=249200 176960 0 180 $X=244850 $Y=171840
X10087 1364 1362 DECAP7JI3V $T=249200 176960 1 0 $X=248770 $Y=171840
X10088 1364 1362 DECAP7JI3V $T=251440 96320 1 0 $X=251010 $Y=91200
X10089 1364 1362 DECAP7JI3V $T=254240 185920 1 0 $X=253810 $Y=180800
X10090 1364 1362 DECAP7JI3V $T=258720 96320 0 0 $X=258290 $Y=95680
X10091 1364 1362 DECAP7JI3V $T=262640 96320 0 0 $X=262210 $Y=95680
X10092 1364 1362 DECAP7JI3V $T=266560 96320 0 0 $X=266130 $Y=95680
X10093 1364 1362 DECAP7JI3V $T=267120 78400 0 0 $X=266690 $Y=77760
X10094 1364 1362 DECAP7JI3V $T=267680 78400 1 0 $X=267250 $Y=73280
X10095 1364 1362 DECAP7JI3V $T=270480 24640 0 0 $X=270050 $Y=24000
X10096 1364 1362 DECAP7JI3V $T=270480 96320 0 0 $X=270050 $Y=95680
X10097 1364 1362 DECAP7JI3V $T=271040 78400 0 0 $X=270610 $Y=77760
X10098 1364 1362 DECAP7JI3V $T=271040 141120 1 0 $X=270610 $Y=136000
X10099 1364 1362 DECAP7JI3V $T=271040 141120 0 0 $X=270610 $Y=140480
X10100 1364 1362 DECAP7JI3V $T=271040 150080 1 0 $X=270610 $Y=144960
X10101 1364 1362 DECAP7JI3V $T=276640 203840 1 0 $X=276210 $Y=198720
X10102 1364 1362 DECAP7JI3V $T=280560 203840 1 0 $X=280130 $Y=198720
X10103 1364 1362 DECAP7JI3V $T=284480 203840 1 0 $X=284050 $Y=198720
X10104 1364 1362 DECAP7JI3V $T=285040 105280 1 0 $X=284610 $Y=100160
X10105 1364 1362 DECAP7JI3V $T=285600 185920 1 0 $X=285170 $Y=180800
X10106 1364 1362 DECAP7JI3V $T=288400 203840 1 0 $X=287970 $Y=198720
X10107 1364 1362 DECAP7JI3V $T=288960 105280 1 0 $X=288530 $Y=100160
X10108 1364 1362 DECAP7JI3V $T=291200 42560 1 0 $X=290770 $Y=37440
X10109 1364 1362 DECAP7JI3V $T=292320 132160 0 0 $X=291890 $Y=131520
X10110 1364 1362 DECAP7JI3V $T=297360 176960 0 0 $X=296930 $Y=176320
X10111 1364 1362 DECAP7JI3V $T=302960 96320 0 0 $X=302530 $Y=95680
X10112 1364 1362 DECAP7JI3V $T=306880 96320 0 0 $X=306450 $Y=95680
X10113 1364 1362 DECAP7JI3V $T=310240 159040 1 0 $X=309810 $Y=153920
X10114 1364 1362 DECAP7JI3V $T=310800 96320 0 0 $X=310370 $Y=95680
X10115 1364 1362 DECAP7JI3V $T=314720 78400 0 0 $X=314290 $Y=77760
X10116 1364 1362 DECAP7JI3V $T=316400 87360 0 0 $X=315970 $Y=86720
X10117 1364 1362 DECAP7JI3V $T=318640 141120 0 0 $X=318210 $Y=140480
X10118 1364 1362 DECAP7JI3V $T=320320 87360 0 0 $X=319890 $Y=86720
X10119 1364 1362 DECAP7JI3V $T=323120 194880 1 0 $X=322690 $Y=189760
X10120 1364 1362 DECAP7JI3V $T=324240 87360 0 0 $X=323810 $Y=86720
X10121 1364 1362 DECAP7JI3V $T=325360 123200 1 0 $X=324930 $Y=118080
X10122 1364 1362 DECAP7JI3V $T=326480 42560 0 0 $X=326050 $Y=41920
X10123 1364 1362 DECAP7JI3V $T=327040 194880 1 0 $X=326610 $Y=189760
X10124 1364 1362 DECAP7JI3V $T=329840 203840 1 0 $X=329410 $Y=198720
X10125 1364 1362 DECAP7JI3V $T=333760 60480 0 0 $X=333330 $Y=59840
X10126 1364 1362 DECAP7JI3V $T=337680 60480 0 0 $X=337250 $Y=59840
X10127 1364 1362 DECAP7JI3V $T=342720 51520 1 0 $X=342290 $Y=46400
X10128 1364 1362 DECAP7JI3V $T=343280 69440 1 0 $X=342850 $Y=64320
X10129 1364 1362 DECAP7JI3V $T=344400 78400 0 0 $X=343970 $Y=77760
X10130 1364 1362 DECAP7JI3V $T=344400 96320 0 0 $X=343970 $Y=95680
X10131 1364 1362 DECAP7JI3V $T=344960 168000 0 0 $X=344530 $Y=167360
X10132 1364 1362 DECAP7JI3V $T=345520 96320 1 0 $X=345090 $Y=91200
X10133 1364 1362 DECAP7JI3V $T=345520 114240 0 0 $X=345090 $Y=113600
X10134 1364 1362 DECAP7JI3V $T=347200 69440 1 0 $X=346770 $Y=64320
X10135 1364 1362 DECAP7JI3V $T=348320 51520 0 0 $X=347890 $Y=50880
X10136 1364 1362 DECAP7JI3V $T=348320 78400 0 0 $X=347890 $Y=77760
X10137 1364 1362 DECAP7JI3V $T=348320 96320 0 0 $X=347890 $Y=95680
X10138 1364 1362 DECAP7JI3V $T=349440 96320 1 0 $X=349010 $Y=91200
X10139 1364 1362 DECAP7JI3V $T=349440 114240 0 0 $X=349010 $Y=113600
X10140 1364 1362 DECAP7JI3V $T=349440 176960 1 0 $X=349010 $Y=171840
X10141 1364 1362 DECAP7JI3V $T=350000 33600 1 0 $X=349570 $Y=28480
X10142 1364 1362 DECAP7JI3V $T=351120 69440 1 0 $X=350690 $Y=64320
X10143 1364 1362 DECAP7JI3V $T=351680 168000 1 0 $X=351250 $Y=162880
X10144 1364 1362 DECAP7JI3V $T=351680 176960 0 0 $X=351250 $Y=176320
X10145 1364 1362 DECAP7JI3V $T=352240 60480 1 0 $X=351810 $Y=55360
X10146 1364 1362 DECAP7JI3V $T=352240 78400 0 0 $X=351810 $Y=77760
X10147 1364 1362 DECAP7JI3V $T=352240 87360 1 0 $X=351810 $Y=82240
X10148 1364 1362 DECAP7JI3V $T=352240 87360 0 0 $X=351810 $Y=86720
X10149 1364 1362 DECAP7JI3V $T=352240 96320 0 0 $X=351810 $Y=95680
X10150 1364 1362 DECAP7JI3V $T=352240 123200 1 0 $X=351810 $Y=118080
X10151 1364 1362 DECAP7JI3V $T=352240 123200 0 0 $X=351810 $Y=122560
X10152 1364 1362 DECAP7JI3V $T=352240 141120 0 0 $X=351810 $Y=140480
X10153 1364 1362 DECAP7JI3V $T=352240 159040 0 0 $X=351810 $Y=158400
X10154 1364 1362 DECAP7JI3V $T=353360 96320 1 0 $X=352930 $Y=91200
X10155 1364 1362 DECAP7JI3V $T=353360 114240 1 0 $X=352930 $Y=109120
X10156 1364 1362 DECAP7JI3V $T=353360 114240 0 0 $X=352930 $Y=113600
X10157 1364 1362 DECAP7JI3V $T=353360 176960 1 0 $X=352930 $Y=171840
X10158 1364 1362 DECAP7JI3V $T=353920 33600 1 0 $X=353490 $Y=28480
X10159 1364 1362 DECAP7JI3V $T=355040 132160 1 0 $X=354610 $Y=127040
X10160 1364 1362 DECAP7JI3V $T=355600 176960 0 0 $X=355170 $Y=176320
X10161 1364 1362 DECAP7JI3V $T=356160 60480 1 0 $X=355730 $Y=55360
X10162 1364 1362 DECAP7JI3V $T=356160 78400 0 0 $X=355730 $Y=77760
X10163 1364 1362 DECAP7JI3V $T=356160 87360 1 0 $X=355730 $Y=82240
X10164 1364 1362 DECAP7JI3V $T=356160 87360 0 0 $X=355730 $Y=86720
X10165 1364 1362 DECAP7JI3V $T=356160 96320 0 0 $X=355730 $Y=95680
X10166 1364 1362 DECAP7JI3V $T=356160 123200 1 0 $X=355730 $Y=118080
X10167 1364 1362 DECAP7JI3V $T=356160 123200 0 0 $X=355730 $Y=122560
X10168 1364 1362 DECAP7JI3V $T=357280 176960 1 0 $X=356850 $Y=171840
X10169 1364 1362 DECAP7JI3V $T=373520 168000 1 0 $X=373090 $Y=162880
X10170 1364 1362 DECAP7JI3V $T=376320 51520 0 0 $X=375890 $Y=50880
X10171 1364 1362 DECAP7JI3V $T=381360 114240 1 0 $X=380930 $Y=109120
X10172 1364 1362 DECAP7JI3V $T=382480 105280 1 0 $X=382050 $Y=100160
X10173 1364 1362 DECAP7JI3V $T=386400 105280 1 0 $X=385970 $Y=100160
X10174 1364 1362 DECAP7JI3V $T=388640 96320 1 0 $X=388210 $Y=91200
X10175 1364 1362 DECAP7JI3V $T=390320 105280 1 0 $X=389890 $Y=100160
X10176 1364 1362 DECAP7JI3V $T=394240 105280 1 0 $X=393810 $Y=100160
X10177 1364 1362 DECAP7JI3V $T=416640 33600 1 0 $X=416210 $Y=28480
X10178 1364 1362 DECAP7JI3V $T=416640 78400 1 0 $X=416210 $Y=73280
X10179 1364 1362 DECAP7JI3V $T=416640 96320 1 0 $X=416210 $Y=91200
X10180 1364 1362 DECAP7JI3V $T=416640 212800 0 0 $X=416210 $Y=212160
X10181 1364 1362 DECAP7JI3V $T=419440 114240 0 0 $X=419010 $Y=113600
X10182 1364 1362 DECAP7JI3V $T=419440 123200 0 0 $X=419010 $Y=122560
X10183 1364 1362 DECAP7JI3V $T=419440 159040 0 0 $X=419010 $Y=158400
X10184 1364 1362 DECAP7JI3V $T=420560 33600 1 0 $X=420130 $Y=28480
X10185 1364 1362 DECAP7JI3V $T=420560 78400 1 0 $X=420130 $Y=73280
X10186 1364 1362 DECAP7JI3V $T=420560 87360 1 0 $X=420130 $Y=82240
X10187 1364 1362 DECAP7JI3V $T=420560 96320 1 0 $X=420130 $Y=91200
X10188 1364 1362 DECAP7JI3V $T=420560 105280 0 0 $X=420130 $Y=104640
X10189 1364 1362 DECAP7JI3V $T=420560 114240 1 0 $X=420130 $Y=109120
X10190 1364 1362 DECAP7JI3V $T=420560 194880 1 0 $X=420130 $Y=189760
X10191 1364 1362 DECAP7JI3V $T=420560 212800 0 0 $X=420130 $Y=212160
X10192 1364 1362 DECAP7JI3V $T=423360 24640 0 0 $X=422930 $Y=24000
X10193 1364 1362 DECAP7JI3V $T=423360 114240 0 0 $X=422930 $Y=113600
X10194 1364 1362 DECAP7JI3V $T=423360 123200 0 0 $X=422930 $Y=122560
X10195 1364 1362 DECAP7JI3V $T=423360 159040 0 0 $X=422930 $Y=158400
X10196 1364 1362 DECAP7JI3V $T=423360 176960 1 0 $X=422930 $Y=171840
X10197 1364 1362 DECAP7JI3V $T=424480 33600 1 0 $X=424050 $Y=28480
X10198 1364 1362 DECAP7JI3V $T=424480 78400 1 0 $X=424050 $Y=73280
X10199 1364 1362 DECAP7JI3V $T=424480 87360 1 0 $X=424050 $Y=82240
X10200 1364 1362 DECAP7JI3V $T=424480 96320 1 0 $X=424050 $Y=91200
X10201 1364 1362 DECAP7JI3V $T=424480 105280 0 0 $X=424050 $Y=104640
X10202 1364 1362 DECAP7JI3V $T=424480 114240 1 0 $X=424050 $Y=109120
X10203 1364 1362 DECAP7JI3V $T=424480 123200 1 0 $X=424050 $Y=118080
X10204 1364 1362 DECAP7JI3V $T=424480 141120 1 0 $X=424050 $Y=136000
X10205 1364 1362 DECAP7JI3V $T=424480 194880 1 0 $X=424050 $Y=189760
X10206 1364 1362 DECAP7JI3V $T=424480 212800 0 0 $X=424050 $Y=212160
X10207 1364 1362 DECAP7JI3V $T=427280 24640 0 0 $X=426850 $Y=24000
X10208 1364 1362 DECAP7JI3V $T=427280 33600 0 0 $X=426850 $Y=32960
X10209 1364 1362 DECAP7JI3V $T=427280 42560 1 0 $X=426850 $Y=37440
X10210 1364 1362 DECAP7JI3V $T=427280 42560 0 0 $X=426850 $Y=41920
X10211 1364 1362 DECAP7JI3V $T=427280 51520 1 0 $X=426850 $Y=46400
X10212 1364 1362 DECAP7JI3V $T=427280 51520 0 0 $X=426850 $Y=50880
X10213 1364 1362 DECAP7JI3V $T=427280 60480 1 0 $X=426850 $Y=55360
X10214 1364 1362 DECAP7JI3V $T=427280 60480 0 0 $X=426850 $Y=59840
X10215 1364 1362 DECAP7JI3V $T=427280 69440 1 0 $X=426850 $Y=64320
X10216 1364 1362 DECAP7JI3V $T=427280 69440 0 0 $X=426850 $Y=68800
X10217 1364 1362 DECAP7JI3V $T=427280 87360 0 0 $X=426850 $Y=86720
X10218 1364 1362 DECAP7JI3V $T=427280 105280 1 0 $X=426850 $Y=100160
X10219 1364 1362 DECAP7JI3V $T=427280 114240 0 0 $X=426850 $Y=113600
X10220 1364 1362 DECAP7JI3V $T=427280 123200 0 0 $X=426850 $Y=122560
X10221 1364 1362 DECAP7JI3V $T=427280 159040 0 0 $X=426850 $Y=158400
X10222 1364 1362 DECAP7JI3V $T=427280 168000 0 0 $X=426850 $Y=167360
X10223 1364 1362 DECAP7JI3V $T=427280 176960 1 0 $X=426850 $Y=171840
X10224 1364 1362 DECAP7JI3V $T=427280 194880 0 0 $X=426850 $Y=194240
X10225 1364 1362 DECAP7JI3V $T=428400 24640 1 0 $X=427970 $Y=19520
X10226 1364 1362 DECAP7JI3V $T=428400 33600 1 0 $X=427970 $Y=28480
X10227 1364 1362 DECAP7JI3V $T=428400 78400 1 0 $X=427970 $Y=73280
X10228 1364 1362 DECAP7JI3V $T=428400 78400 0 0 $X=427970 $Y=77760
X10229 1364 1362 DECAP7JI3V $T=428400 87360 1 0 $X=427970 $Y=82240
X10230 1364 1362 DECAP7JI3V $T=428400 96320 1 0 $X=427970 $Y=91200
X10231 1364 1362 DECAP7JI3V $T=428400 96320 0 0 $X=427970 $Y=95680
X10232 1364 1362 DECAP7JI3V $T=428400 105280 0 0 $X=427970 $Y=104640
X10233 1364 1362 DECAP7JI3V $T=428400 114240 1 0 $X=427970 $Y=109120
X10234 1364 1362 DECAP7JI3V $T=428400 123200 1 0 $X=427970 $Y=118080
X10235 1364 1362 DECAP7JI3V $T=428400 141120 1 0 $X=427970 $Y=136000
X10236 1364 1362 DECAP7JI3V $T=428400 168000 1 0 $X=427970 $Y=162880
X10237 1364 1362 DECAP7JI3V $T=428400 194880 1 0 $X=427970 $Y=189760
X10238 1364 1362 DECAP7JI3V $T=428400 212800 1 0 $X=427970 $Y=207680
X10239 1364 1362 DECAP7JI3V $T=428400 212800 0 0 $X=427970 $Y=212160
X10240 1364 1362 DECAP7JI3V $T=431200 24640 0 0 $X=430770 $Y=24000
X10241 1364 1362 DECAP7JI3V $T=431200 33600 0 0 $X=430770 $Y=32960
X10242 1364 1362 DECAP7JI3V $T=431200 42560 1 0 $X=430770 $Y=37440
X10243 1364 1362 DECAP7JI3V $T=431200 42560 0 0 $X=430770 $Y=41920
X10244 1364 1362 DECAP7JI3V $T=431200 51520 1 0 $X=430770 $Y=46400
X10245 1364 1362 DECAP7JI3V $T=431200 51520 0 0 $X=430770 $Y=50880
X10246 1364 1362 DECAP7JI3V $T=431200 60480 1 0 $X=430770 $Y=55360
X10247 1364 1362 DECAP7JI3V $T=431200 60480 0 0 $X=430770 $Y=59840
X10248 1364 1362 DECAP7JI3V $T=431200 69440 1 0 $X=430770 $Y=64320
X10249 1364 1362 DECAP7JI3V $T=431200 69440 0 0 $X=430770 $Y=68800
X10250 1364 1362 DECAP7JI3V $T=431200 87360 0 0 $X=430770 $Y=86720
X10251 1364 1362 DECAP7JI3V $T=431200 105280 1 0 $X=430770 $Y=100160
X10252 1364 1362 DECAP7JI3V $T=431200 114240 0 0 $X=430770 $Y=113600
X10253 1364 1362 DECAP7JI3V $T=431200 123200 0 0 $X=430770 $Y=122560
X10254 1364 1362 DECAP7JI3V $T=431200 150080 0 0 $X=430770 $Y=149440
X10255 1364 1362 DECAP7JI3V $T=431200 159040 0 0 $X=430770 $Y=158400
X10256 1364 1362 DECAP7JI3V $T=431200 168000 0 0 $X=430770 $Y=167360
X10257 1364 1362 DECAP7JI3V $T=431200 176960 1 0 $X=430770 $Y=171840
X10258 1364 1362 DECAP7JI3V $T=431200 176960 0 0 $X=430770 $Y=176320
X10259 1364 1362 DECAP7JI3V $T=431200 185920 1 0 $X=430770 $Y=180800
X10260 1364 1362 DECAP7JI3V $T=431200 194880 0 0 $X=430770 $Y=194240
X10261 1364 1362 DECAP7JI3V $T=431200 203840 1 0 $X=430770 $Y=198720
X10262 1364 1362 DECAP5JI3V $T=20160 105280 0 0 $X=19730 $Y=104640
X10263 1364 1362 DECAP5JI3V $T=20160 114240 1 0 $X=19730 $Y=109120
X10264 1364 1362 DECAP5JI3V $T=20160 123200 0 0 $X=19730 $Y=122560
X10265 1364 1362 DECAP5JI3V $T=20160 132160 1 0 $X=19730 $Y=127040
X10266 1364 1362 DECAP5JI3V $T=20160 132160 0 0 $X=19730 $Y=131520
X10267 1364 1362 DECAP5JI3V $T=20160 194880 1 0 $X=19730 $Y=189760
X10268 1364 1362 DECAP5JI3V $T=36960 114240 0 0 $X=36530 $Y=113600
X10269 1364 1362 DECAP5JI3V $T=42000 42560 1 0 $X=41570 $Y=37440
X10270 1364 1362 DECAP5JI3V $T=42000 42560 0 0 $X=41570 $Y=41920
X10271 1364 1362 DECAP5JI3V $T=42000 51520 1 0 $X=41570 $Y=46400
X10272 1364 1362 DECAP5JI3V $T=42000 51520 0 0 $X=41570 $Y=50880
X10273 1364 1362 DECAP5JI3V $T=42560 60480 1 0 $X=42130 $Y=55360
X10274 1364 1362 DECAP5JI3V $T=48160 176960 1 0 $X=47730 $Y=171840
X10275 1364 1362 DECAP5JI3V $T=48160 203840 1 0 $X=47730 $Y=198720
X10276 1364 1362 DECAP5JI3V $T=54320 24640 1 0 $X=53890 $Y=19520
X10277 1364 1362 DECAP5JI3V $T=59920 42560 1 0 $X=59490 $Y=37440
X10278 1364 1362 DECAP5JI3V $T=60480 60480 0 0 $X=60050 $Y=59840
X10279 1364 1362 DECAP5JI3V $T=62160 78400 0 0 $X=61730 $Y=77760
X10280 1364 1362 DECAP5JI3V $T=62160 87360 0 0 $X=61730 $Y=86720
X10281 1364 1362 DECAP5JI3V $T=62720 105280 0 0 $X=62290 $Y=104640
X10282 1364 1362 DECAP5JI3V $T=63280 114240 0 0 $X=62850 $Y=113600
X10283 1364 1362 DECAP5JI3V $T=67760 159040 1 0 $X=67330 $Y=153920
X10284 1364 1362 DECAP5JI3V $T=72240 212800 1 0 $X=71810 $Y=207680
X10285 1364 1362 DECAP5JI3V $T=94080 51520 1 0 $X=93650 $Y=46400
X10286 1364 1362 DECAP5JI3V $T=94080 51520 0 0 $X=93650 $Y=50880
X10287 1364 1362 DECAP5JI3V $T=94080 60480 1 0 $X=93650 $Y=55360
X10288 1364 1362 DECAP5JI3V $T=95760 150080 1 0 $X=95330 $Y=144960
X10289 1364 1362 DECAP5JI3V $T=98560 185920 1 0 $X=98130 $Y=180800
X10290 1364 1362 DECAP5JI3V $T=100240 105280 1 0 $X=99810 $Y=100160
X10291 1364 1362 DECAP5JI3V $T=100240 123200 0 0 $X=99810 $Y=122560
X10292 1364 1362 DECAP5JI3V $T=100240 132160 1 0 $X=99810 $Y=127040
X10293 1364 1362 DECAP5JI3V $T=100240 141120 0 0 $X=99810 $Y=140480
X10294 1364 1362 DECAP5JI3V $T=100240 159040 1 0 $X=99810 $Y=153920
X10295 1364 1362 DECAP5JI3V $T=107520 105280 0 0 $X=107090 $Y=104640
X10296 1364 1362 DECAP5JI3V $T=108080 87360 0 0 $X=107650 $Y=86720
X10297 1364 1362 DECAP5JI3V $T=108640 78400 0 0 $X=108210 $Y=77760
X10298 1364 1362 DECAP5JI3V $T=110880 114240 1 0 $X=110450 $Y=109120
X10299 1364 1362 DECAP5JI3V $T=115360 114240 0 0 $X=114930 $Y=113600
X10300 1364 1362 DECAP5JI3V $T=121520 24640 1 180 $X=118290 $Y=24000
X10301 1364 1362 DECAP5JI3V $T=119280 168000 0 0 $X=118850 $Y=167360
X10302 1364 1362 DECAP5JI3V $T=134960 24640 1 0 $X=134530 $Y=19520
X10303 1364 1362 DECAP5JI3V $T=140000 78400 0 0 $X=139570 $Y=77760
X10304 1364 1362 DECAP5JI3V $T=140000 87360 0 0 $X=139570 $Y=86720
X10305 1364 1362 DECAP5JI3V $T=142800 69440 0 0 $X=142370 $Y=68800
X10306 1364 1362 DECAP5JI3V $T=156240 212800 0 0 $X=155810 $Y=212160
X10307 1364 1362 DECAP5JI3V $T=159600 78400 1 0 $X=159170 $Y=73280
X10308 1364 1362 DECAP5JI3V $T=163520 168000 1 0 $X=163090 $Y=162880
X10309 1364 1362 DECAP5JI3V $T=166320 33600 0 0 $X=165890 $Y=32960
X10310 1364 1362 DECAP5JI3V $T=179760 60480 1 0 $X=179330 $Y=55360
X10311 1364 1362 DECAP5JI3V $T=181440 168000 1 0 $X=181010 $Y=162880
X10312 1364 1362 DECAP5JI3V $T=184240 87360 1 0 $X=183810 $Y=82240
X10313 1364 1362 DECAP5JI3V $T=184800 42560 1 0 $X=184370 $Y=37440
X10314 1364 1362 DECAP5JI3V $T=185360 132160 1 0 $X=184930 $Y=127040
X10315 1364 1362 DECAP5JI3V $T=188720 212800 1 0 $X=188290 $Y=207680
X10316 1364 1362 DECAP5JI3V $T=197680 51520 1 0 $X=197250 $Y=46400
X10317 1364 1362 DECAP5JI3V $T=197680 51520 0 0 $X=197250 $Y=50880
X10318 1364 1362 DECAP5JI3V $T=224000 51520 1 0 $X=223570 $Y=46400
X10319 1364 1362 DECAP5JI3V $T=224000 60480 0 0 $X=223570 $Y=59840
X10320 1364 1362 DECAP5JI3V $T=224000 176960 0 0 $X=223570 $Y=176320
X10321 1364 1362 DECAP5JI3V $T=224000 185920 1 0 $X=223570 $Y=180800
X10322 1364 1362 DECAP5JI3V $T=228480 141120 0 0 $X=228050 $Y=140480
X10323 1364 1362 DECAP5JI3V $T=228480 150080 0 0 $X=228050 $Y=149440
X10324 1364 1362 DECAP5JI3V $T=229040 33600 1 0 $X=228610 $Y=28480
X10325 1364 1362 DECAP5JI3V $T=229040 212800 0 0 $X=228610 $Y=212160
X10326 1364 1362 DECAP5JI3V $T=230160 24640 0 0 $X=229730 $Y=24000
X10327 1364 1362 DECAP5JI3V $T=230160 87360 1 0 $X=229730 $Y=82240
X10328 1364 1362 DECAP5JI3V $T=230720 168000 0 0 $X=230290 $Y=167360
X10329 1364 1362 DECAP5JI3V $T=231840 114240 1 0 $X=231410 $Y=109120
X10330 1364 1362 DECAP5JI3V $T=237440 123200 0 0 $X=237010 $Y=122560
X10331 1364 1362 DECAP5JI3V $T=244160 33600 1 0 $X=243730 $Y=28480
X10332 1364 1362 DECAP5JI3V $T=251440 114240 1 0 $X=251010 $Y=109120
X10333 1364 1362 DECAP5JI3V $T=263760 176960 1 0 $X=263330 $Y=171840
X10334 1364 1362 DECAP5JI3V $T=272160 132160 1 0 $X=271730 $Y=127040
X10335 1364 1362 DECAP5JI3V $T=273280 60480 1 0 $X=272850 $Y=55360
X10336 1364 1362 DECAP5JI3V $T=274400 123200 0 0 $X=273970 $Y=122560
X10337 1364 1362 DECAP5JI3V $T=276080 203840 0 0 $X=275650 $Y=203200
X10338 1364 1362 DECAP5JI3V $T=277760 132160 0 0 $X=277330 $Y=131520
X10339 1364 1362 DECAP5JI3V $T=278320 33600 0 0 $X=277890 $Y=32960
X10340 1364 1362 DECAP5JI3V $T=285040 33600 1 0 $X=284610 $Y=28480
X10341 1364 1362 DECAP5JI3V $T=285600 114240 0 0 $X=285170 $Y=113600
X10342 1364 1362 DECAP5JI3V $T=294000 51520 0 180 $X=290770 $Y=46400
X10343 1364 1362 DECAP5JI3V $T=291200 51520 0 0 $X=290770 $Y=50880
X10344 1364 1362 DECAP5JI3V $T=291200 60480 1 0 $X=290770 $Y=55360
X10345 1364 1362 DECAP5JI3V $T=291200 60480 0 0 $X=290770 $Y=59840
X10346 1364 1362 DECAP5JI3V $T=291760 96320 1 0 $X=291330 $Y=91200
X10347 1364 1362 DECAP5JI3V $T=299040 159040 1 0 $X=298610 $Y=153920
X10348 1364 1362 DECAP5JI3V $T=301840 33600 0 0 $X=301410 $Y=32960
X10349 1364 1362 DECAP5JI3V $T=306880 194880 1 0 $X=306450 $Y=189760
X10350 1364 1362 DECAP5JI3V $T=309120 60480 0 0 $X=308690 $Y=59840
X10351 1364 1362 DECAP5JI3V $T=312480 212800 1 0 $X=312050 $Y=207680
X10352 1364 1362 DECAP5JI3V $T=314160 114240 0 0 $X=313730 $Y=113600
X10353 1364 1362 DECAP5JI3V $T=317520 24640 0 0 $X=317090 $Y=24000
X10354 1364 1362 DECAP5JI3V $T=327040 78400 1 0 $X=326610 $Y=73280
X10355 1364 1362 DECAP5JI3V $T=327040 194880 0 0 $X=326610 $Y=194240
X10356 1364 1362 DECAP5JI3V $T=328720 69440 0 0 $X=328290 $Y=68800
X10357 1364 1362 DECAP5JI3V $T=342720 212800 1 0 $X=342290 $Y=207680
X10358 1364 1362 DECAP5JI3V $T=352240 51520 0 0 $X=351810 $Y=50880
X10359 1364 1362 DECAP5JI3V $T=355040 159040 1 0 $X=354610 $Y=153920
X10360 1364 1362 DECAP5JI3V $T=355600 141120 1 0 $X=355170 $Y=136000
X10361 1364 1362 DECAP5JI3V $T=355600 150080 1 0 $X=355170 $Y=144960
X10362 1364 1362 DECAP5JI3V $T=355600 168000 1 0 $X=355170 $Y=162880
X10363 1364 1362 DECAP5JI3V $T=357280 96320 1 0 $X=356850 $Y=91200
X10364 1364 1362 DECAP5JI3V $T=357280 114240 0 0 $X=356850 $Y=113600
X10365 1364 1362 DECAP5JI3V $T=357840 33600 1 0 $X=357410 $Y=28480
X10366 1364 1362 DECAP5JI3V $T=358400 105280 1 0 $X=357970 $Y=100160
X10367 1364 1362 DECAP5JI3V $T=362880 51520 0 180 $X=359650 $Y=46400
X10368 1364 1362 DECAP5JI3V $T=360080 60480 1 0 $X=359650 $Y=55360
X10369 1364 1362 DECAP5JI3V $T=377440 60480 0 0 $X=377010 $Y=59840
X10370 1364 1362 DECAP5JI3V $T=383040 132160 0 180 $X=379810 $Y=127040
X10371 1364 1362 DECAP5JI3V $T=381360 105280 0 0 $X=380930 $Y=104640
X10372 1364 1362 DECAP5JI3V $T=381360 123200 1 0 $X=380930 $Y=118080
X10373 1364 1362 DECAP5JI3V $T=381920 114240 0 0 $X=381490 $Y=113600
X10374 1364 1362 DECAP5JI3V $T=381920 141120 0 0 $X=381490 $Y=140480
X10375 1364 1362 DECAP5JI3V $T=385840 33600 1 0 $X=385410 $Y=28480
X10376 1364 1362 DECAP5JI3V $T=393680 150080 1 180 $X=390450 $Y=149440
X10377 1364 1362 DECAP5JI3V $T=392560 96320 1 0 $X=392130 $Y=91200
X10378 1364 1362 DECAP5JI3V $T=395360 42560 1 0 $X=394930 $Y=37440
X10379 1364 1362 DECAP5JI3V $T=395360 42560 0 0 $X=394930 $Y=41920
X10380 1364 1362 DECAP5JI3V $T=395360 60480 1 0 $X=394930 $Y=55360
X10381 1364 1362 DECAP5JI3V $T=395360 60480 0 0 $X=394930 $Y=59840
X10382 1364 1362 DECAP5JI3V $T=395360 69440 1 0 $X=394930 $Y=64320
X10383 1364 1362 DECAP5JI3V $T=395360 69440 0 0 $X=394930 $Y=68800
X10384 1364 1362 DECAP5JI3V $T=409360 24640 1 180 $X=406130 $Y=24000
X10385 1364 1362 DECAP5JI3V $T=432320 24640 1 0 $X=431890 $Y=19520
X10386 1364 1362 DECAP5JI3V $T=432320 33600 1 0 $X=431890 $Y=28480
X10387 1364 1362 DECAP5JI3V $T=432320 78400 1 0 $X=431890 $Y=73280
X10388 1364 1362 DECAP5JI3V $T=432320 78400 0 0 $X=431890 $Y=77760
X10389 1364 1362 DECAP5JI3V $T=432320 87360 1 0 $X=431890 $Y=82240
X10390 1364 1362 DECAP5JI3V $T=432320 96320 1 0 $X=431890 $Y=91200
X10391 1364 1362 DECAP5JI3V $T=432320 96320 0 0 $X=431890 $Y=95680
X10392 1364 1362 DECAP5JI3V $T=432320 105280 0 0 $X=431890 $Y=104640
X10393 1364 1362 DECAP5JI3V $T=432320 114240 1 0 $X=431890 $Y=109120
X10394 1364 1362 DECAP5JI3V $T=432320 123200 1 0 $X=431890 $Y=118080
X10395 1364 1362 DECAP5JI3V $T=432320 132160 1 0 $X=431890 $Y=127040
X10396 1364 1362 DECAP5JI3V $T=432320 141120 1 0 $X=431890 $Y=136000
X10397 1364 1362 DECAP5JI3V $T=432320 159040 1 0 $X=431890 $Y=153920
X10398 1364 1362 DECAP5JI3V $T=432320 168000 1 0 $X=431890 $Y=162880
X10399 1364 1362 DECAP5JI3V $T=432320 194880 1 0 $X=431890 $Y=189760
X10400 1364 1362 DECAP5JI3V $T=432320 212800 1 0 $X=431890 $Y=207680
X10401 1364 1362 DECAP5JI3V $T=432320 212800 0 0 $X=431890 $Y=212160
X10402 1364 1362 DECAP10JI3V $T=20160 114240 0 0 $X=19730 $Y=113600
X10403 1364 1362 DECAP10JI3V $T=20160 123200 1 0 $X=19730 $Y=118080
X10404 1364 1362 DECAP10JI3V $T=20160 159040 1 0 $X=19730 $Y=153920
X10405 1364 1362 DECAP10JI3V $T=20160 176960 0 0 $X=19730 $Y=176320
X10406 1364 1362 DECAP10JI3V $T=20160 185920 0 0 $X=19730 $Y=185280
X10407 1364 1362 DECAP10JI3V $T=34160 24640 0 0 $X=33730 $Y=24000
X10408 1364 1362 DECAP10JI3V $T=34160 87360 1 0 $X=33730 $Y=82240
X10409 1364 1362 DECAP10JI3V $T=34160 194880 0 0 $X=33730 $Y=194240
X10410 1364 1362 DECAP10JI3V $T=39760 123200 0 0 $X=39330 $Y=122560
X10411 1364 1362 DECAP10JI3V $T=76160 203840 1 0 $X=75730 $Y=198720
X10412 1364 1362 DECAP10JI3V $T=77840 141120 0 0 $X=77410 $Y=140480
X10413 1364 1362 DECAP10JI3V $T=90720 176960 1 0 $X=90290 $Y=171840
X10414 1364 1362 DECAP10JI3V $T=92960 168000 0 0 $X=92530 $Y=167360
X10415 1364 1362 DECAP10JI3V $T=95200 159040 0 0 $X=94770 $Y=158400
X10416 1364 1362 DECAP10JI3V $T=95760 176960 0 0 $X=95330 $Y=176320
X10417 1364 1362 DECAP10JI3V $T=100240 194880 1 0 $X=99810 $Y=189760
X10418 1364 1362 DECAP10JI3V $T=140560 176960 1 0 $X=140130 $Y=171840
X10419 1364 1362 DECAP10JI3V $T=151760 132160 0 0 $X=151330 $Y=131520
X10420 1364 1362 DECAP10JI3V $T=152880 87360 1 0 $X=152450 $Y=82240
X10421 1364 1362 DECAP10JI3V $T=204400 123200 1 0 $X=203970 $Y=118080
X10422 1364 1362 DECAP10JI3V $T=212240 42560 1 0 $X=211810 $Y=37440
X10423 1364 1362 DECAP10JI3V $T=221200 51520 0 0 $X=220770 $Y=50880
X10424 1364 1362 DECAP10JI3V $T=223440 78400 0 0 $X=223010 $Y=77760
X10425 1364 1362 DECAP10JI3V $T=223440 87360 0 0 $X=223010 $Y=86720
X10426 1364 1362 DECAP10JI3V $T=223440 96320 0 0 $X=223010 $Y=95680
X10427 1364 1362 DECAP10JI3V $T=223440 105280 0 0 $X=223010 $Y=104640
X10428 1364 1362 DECAP10JI3V $T=223440 132160 0 0 $X=223010 $Y=131520
X10429 1364 1362 DECAP10JI3V $T=223440 159040 1 0 $X=223010 $Y=153920
X10430 1364 1362 DECAP10JI3V $T=224560 176960 1 0 $X=224130 $Y=171840
X10431 1364 1362 DECAP10JI3V $T=226240 123200 1 0 $X=225810 $Y=118080
X10432 1364 1362 DECAP10JI3V $T=228480 141120 1 0 $X=228050 $Y=136000
X10433 1364 1362 DECAP10JI3V $T=243040 150080 1 0 $X=242610 $Y=144960
X10434 1364 1362 DECAP10JI3V $T=245840 96320 1 0 $X=245410 $Y=91200
X10435 1364 1362 DECAP10JI3V $T=253120 105280 0 0 $X=252690 $Y=104640
X10436 1364 1362 DECAP10JI3V $T=283360 150080 0 0 $X=282930 $Y=149440
X10437 1364 1362 DECAP10JI3V $T=285600 42560 1 0 $X=285170 $Y=37440
X10438 1364 1362 DECAP10JI3V $T=308560 176960 0 0 $X=308130 $Y=176320
X10439 1364 1362 DECAP10JI3V $T=309120 78400 0 0 $X=308690 $Y=77760
X10440 1364 1362 DECAP10JI3V $T=318640 123200 1 0 $X=318210 $Y=118080
X10441 1364 1362 DECAP10JI3V $T=326480 105280 0 0 $X=326050 $Y=104640
X10442 1364 1362 DECAP10JI3V $T=338800 78400 0 0 $X=338370 $Y=77760
X10443 1364 1362 DECAP10JI3V $T=340480 33600 1 0 $X=340050 $Y=28480
X10444 1364 1362 DECAP10JI3V $T=347760 114240 1 0 $X=347330 $Y=109120
X10445 1364 1362 DECAP10JI3V $T=352240 42560 1 0 $X=351810 $Y=37440
X10446 1364 1362 DECAP10JI3V $T=352240 105280 0 0 $X=351810 $Y=104640
X10447 1364 1362 DECAP10JI3V $T=352240 185920 0 0 $X=351810 $Y=185280
X10448 1364 1362 DECAP10JI3V $T=352800 168000 0 0 $X=352370 $Y=167360
X10449 1364 1362 DECAP10JI3V $T=356720 42560 0 0 $X=356290 $Y=41920
X10450 1364 1362 DECAP10JI3V $T=356720 60480 0 0 $X=356290 $Y=59840
X10451 1364 1362 DECAP10JI3V $T=373520 185920 0 180 $X=367490 $Y=180800
X10452 1364 1362 DECAP10JI3V $T=371280 69440 1 0 $X=370850 $Y=64320
X10453 1364 1362 DECAP10JI3V $T=413840 123200 0 0 $X=413410 $Y=122560
X10454 1364 1362 DECAP10JI3V $T=413840 159040 0 0 $X=413410 $Y=158400
X10455 1364 1362 DECAP10JI3V $T=421680 33600 0 0 $X=421250 $Y=32960
X10456 1364 1362 DECAP10JI3V $T=421680 60480 1 0 $X=421250 $Y=55360
X10457 1364 1362 DECAP10JI3V $T=421680 87360 0 0 $X=421250 $Y=86720
X10458 1364 1362 DECAP10JI3V $T=421680 168000 0 0 $X=421250 $Y=167360
D0 1363 1364 p_ddnwmv AREA=8.49716e-08 PJ=0.00124444 perimeter=0.00124444 $X=17730 $Y=17520 $dt=2
D1 1362 1364 p_dipdnwmv AREA=1.68269e-09 PJ=0.000846738 perimeter=0.000846738 $X=24380 $Y=192640 $dt=3
D2 1362 1364 p_dipdnwmv AREA=1.71436e-09 PJ=0.000856626 perimeter=0.000856626 $X=29010 $Y=138870 $dt=3
D3 1362 1364 p_dipdnwmv AREA=1.70244e-09 PJ=0.00085168 perimeter=0.00085168 $X=30130 $Y=120950 $dt=3
D4 1362 1364 p_dipdnwmv AREA=1.7101e-09 PJ=0.000852491 perimeter=0.000852491 $X=46940 $Y=94080 $dt=3
D5 1362 1364 p_dipdnwmv AREA=1.72326e-09 PJ=0.000856437 perimeter=0.000856437 $X=69890 $Y=67190 $dt=3
D6 1362 1364 p_dipdnwmv AREA=1.68194e-09 PJ=0.000847719 perimeter=0.000847719 $X=76460 $Y=210560 $dt=3
D7 1362 1364 p_dipdnwmv AREA=1.72011e-09 PJ=0.000854508 perimeter=0.000854508 $X=85570 $Y=85110 $dt=3
D8 1362 1364 p_dipdnwmv AREA=1.68085e-09 PJ=0.000847368 perimeter=0.000847368 $X=85570 $Y=201590 $dt=3
D9 1362 1364 p_dipdnwmv AREA=1.67889e-09 PJ=0.000849321 perimeter=0.000849321 $X=87810 $Y=165750 $dt=3
D10 1362 1364 p_dipdnwmv AREA=1.7123e-09 PJ=0.000855368 perimeter=0.000855368 $X=89490 $Y=147830 $dt=3
D11 1362 1364 p_dipdnwmv AREA=1.66499e-09 PJ=0.000851237 perimeter=0.000851237 $X=117490 $Y=31350 $dt=3
D12 1362 1364 p_dipdnwmv AREA=1.71216e-09 PJ=0.000861885 perimeter=0.000861885 $X=129810 $Y=40310 $dt=3
D13 1362 1364 p_dipdnwmv AREA=1.67656e-09 PJ=0.000846569 perimeter=0.000846569 $X=132610 $Y=183670 $dt=3
D14 1362 1364 p_dipdnwmv AREA=1.72262e-09 PJ=0.000856557 perimeter=0.000856557 $X=146610 $Y=58230 $dt=3
D15 1362 1364 p_dipdnwmv AREA=1.70024e-09 PJ=0.000851249 perimeter=0.000851249 $X=167890 $Y=111990 $dt=3
D16 1362 1364 p_dipdnwmv AREA=1.71539e-09 PJ=0.000856066 perimeter=0.000856066 $X=175170 $Y=129910 $dt=3
D17 1362 1364 p_dipdnwmv AREA=1.71256e-09 PJ=0.000853309 perimeter=0.000853309 $X=191410 $Y=103030 $dt=3
D18 1362 1364 p_dipdnwmv AREA=1.69697e-09 PJ=0.000852039 perimeter=0.000852039 $X=293890 $Y=156790 $dt=3
D19 1362 1364 p_dipdnwmv AREA=1.67952e-09 PJ=0.000847075 perimeter=0.000847075 $X=344380 $Y=174710 $dt=3
D20 1362 1364 p_dipdnwmv AREA=1.64744e-09 PJ=0.0008401 perimeter=0.0008401 $X=386290 $Y=22390 $dt=3
D21 1362 1364 p_dipdnwmv AREA=1.71423e-09 PJ=0.000853703 perimeter=0.000853703 $X=390210 $Y=76150 $dt=3
D22 1362 1364 p_dipdnwmv AREA=1.72604e-09 PJ=0.000856428 perimeter=0.000856428 $X=413730 $Y=49270 $dt=3
.ends aska_dig
