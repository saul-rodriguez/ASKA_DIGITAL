* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : aska_dig                                     *
* Netlisted  : Mon Jul 15 19:33:54 2024                     *
* PVS Version: 23.10-p043 Mon Oct 2 18:09:08 PDT 2023      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(ne3i) nemi ndiff(D) p1trm(G) ndiff(S) pwitrm(B)
*.DEVTMPLT 1 MP(pe3i) pemi pdiff(D) p1trm(G) pdiff(S) dnwtrm(B)
*.DEVTMPLT 2 D(p_ddnwmv) p_ddnwmv bulk(POS) dnwtrm(NEG)
*.DEVTMPLT 3 D(p_dipdnwmv) p_dipwmv pwitrm(POS) dnwtrm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX2                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX2 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=6
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=6e-07 AD=2.96727e-13 AS=2.88e-13 PD=1.69091e-06 PS=2.16e-06 $X=620 $Y=950 $dt=0
M1 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=7.2e-07 AD=2.016e-13 AS=3.56073e-13 PD=1.512e-06 PS=2.02909e-06 $X=1590 $Y=830 $dt=0
M2 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=4.648e-13 AS=1.344e-13 PD=3.52e-06 PS=1.008e-06 $X=2480 $Y=1070 $dt=0
M3 vdd3i! A 6 vdd3i! pe3i L=3e-07 W=1.1e-06 AD=5.39943e-13 AS=5.28e-13 PD=2.20442e-06 PS=3.16e-06 $X=620 $Y=2410 $dt=1
M4 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=7.16507e-13 PD=1.87971e-06 PS=2.92528e-06 $X=1640 $Y=2410 $dt=1
M5 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=8.6265e-13 AS=2.751e-13 PD=4.56971e-06 PS=1.87971e-06 $X=2480 $Y=2410 $dt=1
.ends BUJI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND2JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND2JI3VX1 vdd3i! gnd3i! A B Q
*.DEVICECLIMB
** N=8 EP=5 FDC=6
M0 7 A 8 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=2.688e-13 PD=8.1e-07 PS=2.08e-06 $X=820 $Y=990 $dt=0
M1 gnd3i! B 7 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=2.57137e-13 AS=7e-14 PD=1.43669e-06 PS=8.1e-07 $X=1420 $Y=990 $dt=0
M2 Q 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=4.08663e-13 PD=2.74e-06 PS=2.28331e-06 $X=2390 $Y=660 $dt=0
M3 8 A vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=7.276e-13 PD=1.24e-06 PS=4.56e-06 $X=580 $Y=2410 $dt=1
M4 vdd3i! B 8 vdd3i! pe3i L=3e-07 W=7e-07 AD=3.64829e-13 AS=1.89e-13 PD=1.6455e-06 PS=1.24e-06 $X=1420 $Y=2410 $dt=1
M5 Q 8 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=7.34871e-13 PD=3.78e-06 PS=3.3145e-06 $X=2440 $Y=2410 $dt=1
.ends AND2JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: EN2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt EN2JI3VX0 vdd3i! gnd3i! A B Q
*.DEVICECLIMB
** N=10 EP=5 FDC=10
M0 8 A 9 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=620 $Y=980 $dt=0
M1 gnd3i! B 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=1220 $Y=980 $dt=0
M2 7 A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=1.134e-13 PD=9.6e-07 PS=9.6e-07 $X=2110 $Y=980 $dt=0
M3 gnd3i! B 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.698e-13 AS=1.134e-13 PD=3.22e-06 PS=9.6e-07 $X=3000 $Y=980 $dt=0
M4 Q 9 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=2.058e-13 PD=1.8e-06 PS=1.82e-06 $X=4440 $Y=1020 $dt=0
M5 9 A vdd3i! vdd3i! pe3i L=3e-07 W=9e-07 AD=3.195e-13 AS=8.517e-13 PD=1.61e-06 PS=4.61e-06 $X=685 $Y=2410 $dt=1
M6 vdd3i! B 9 vdd3i! pe3i L=3e-07 W=9e-07 AD=4.30855e-13 AS=3.195e-13 PD=1.83273e-06 PS=1.61e-06 $X=1695 $Y=2410 $dt=1
M7 10 A vdd3i! vdd3i! pe3i L=3e-07 W=1.3e-06 AD=1.95e-13 AS=6.22345e-13 PD=1.6e-06 PS=2.64727e-06 $X=2825 $Y=2520 $dt=1
M8 Q B 10 vdd3i! pe3i L=3e-07 W=1.3e-06 AD=6.21324e-13 AS=1.95e-13 PD=2.52941e-06 PS=1.6e-06 $X=3425 $Y=2520 $dt=1
M9 vdd3i! 9 Q vdd3i! pe3i L=3e-07 W=9.1e-07 AD=8.0675e-13 AS=4.34926e-13 PD=4.39e-06 PS=1.77059e-06 $X=4575 $Y=2520 $dt=1
.ends EN2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA2I1JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA2I1JI3VX1 vdd3i! gnd3i! AN Q B
*.DEVICECLIMB
** N=8 EP=5 FDC=6
M0 gnd3i! AN 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.44754e-13 AS=2.016e-13 PD=1.25038e-06 PS=1.8e-06 $X=620 $Y=660 $dt=0
M1 7 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=5.18646e-13 PD=1.14e-06 PS=2.64962e-06 $X=1680 $Y=660 $dt=0
M2 Q B 7 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=1.1125e-13 PD=2.74e-06 PS=1.14e-06 $X=2280 $Y=660 $dt=0
M3 vdd3i! AN 8 vdd3i! pe3i L=3e-07 W=7e-07 AD=6.84341e-13 AS=3.36e-13 PD=3.08e-06 PS=2.36e-06 $X=620 $Y=2410 $dt=1
M4 Q 8 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.7e-13 AS=9.7763e-13 PD=1.54e-06 PS=4.4e-06 $X=1510 $Y=2410 $dt=1
M5 vdd3i! B Q vdd3i! pe3i L=3e-07 W=1e-06 AD=9.7763e-13 AS=2.7e-13 PD=4.4e-06 PS=1.54e-06 $X=2350 $Y=2410 $dt=1
.ends NA2I1JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO3I2JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO3I2JI3VX1 vdd3i! gnd3i! AN BN C Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 8 AN 9 gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=6e-14 AS=2.304e-13 PD=7.3e-07 PS=1.92e-06 $X=620 $Y=1070 $dt=0
M1 gnd3i! BN 8 gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=1.98937e-13 AS=6e-14 PD=1.31617e-06 PS=7.3e-07 $X=1220 $Y=1070 $dt=0
M2 Q C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.68863e-13 PD=1.43e-06 PS=2.4404e-06 $X=2060 $Y=660 $dt=0
M3 gnd3i! 9 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.329e-13 AS=2.403e-13 PD=2.77e-06 PS=1.43e-06 $X=2950 $Y=660 $dt=0
M4 9 AN vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=5.71409e-13 PD=1.24e-06 PS=2.5758e-06 $X=560 $Y=2590 $dt=1
M5 vdd3i! BN 9 vdd3i! pe3i L=3e-07 W=7e-07 AD=5.71409e-13 AS=1.89e-13 PD=2.5758e-06 PS=1.24e-06 $X=1400 $Y=2590 $dt=1
M6 10 C vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=1.15098e-12 PD=1.66e-06 PS=5.1884e-06 $X=2330 $Y=2410 $dt=1
M7 Q 9 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=8.46e-13 AS=1.7625e-13 PD=4.02e-06 PS=1.66e-06 $X=2880 $Y=2410 $dt=1
.ends NO3I2JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA2JI3VX1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA2JI3VX1 vdd3i! gnd3i! B Q A
*.DEVICECLIMB
** N=7 EP=5 FDC=4
M0 7 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=6.222e-13 PD=1.14e-06 PS=3.54e-06 $X=670 $Y=660 $dt=0
M1 Q A 7 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=1.1125e-13 PD=2.74e-06 PS=1.14e-06 $X=1270 $Y=660 $dt=0
M2 Q B vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.7e-13 AS=9.404e-13 PD=1.54e-06 PS=5.24e-06 $X=550 $Y=2410 $dt=1
M3 vdd3i! A Q vdd3i! pe3i L=3e-07 W=1e-06 AD=9.404e-13 AS=2.7e-13 PD=5.24e-06 PS=1.54e-06 $X=1390 $Y=2410 $dt=1
.ends NA2JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX1 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=4
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.44533e-13 AS=2.016e-13 PD=1.44667e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=6.6e-07 AD=2.88e-13 AS=3.84267e-13 PD=2.28e-06 PS=2.27333e-06 $X=1590 $Y=890 $dt=0
M2 vdd3i! A 6 vdd3i! pe3i L=3e-07 W=9e-07 AD=4.7931e-13 AS=4.32e-13 PD=1.95649e-06 PS=2.76e-06 $X=620 $Y=2410 $dt=1
M3 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=5.712e-13 AS=7.7739e-13 PD=3.70971e-06 PS=3.17322e-06 $X=1640 $Y=2410 $dt=1
.ends BUJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DFRRQJI3VX4                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DFRRQJI3VX4 vdd3i! gnd3i! RN D C Q
*.DEVICECLIMB
** N=23 EP=6 FDC=36
M0 gnd3i! 17 19 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=4.272e-13 PD=1.43e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 10 RN gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.28952e-13 AS=2.403e-13 PD=2.36956e-06 PS=1.43e-06 $X=1510 $Y=660 $dt=0
M2 18 19 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.55236e-13 PD=6.7e-07 PS=1.11822e-06 $X=2340 $Y=1390 $dt=0
M3 17 9 18 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=2940 $Y=1390 $dt=0
M4 16 15 17 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=3830 $Y=1390 $dt=0
M5 10 D 16 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.835e-13 AS=5.25e-14 PD=2.19e-06 PS=6.7e-07 $X=4430 $Y=1390 $dt=0
M6 gnd3i! C 15 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.659e-13 AS=2.016e-13 PD=1.21e-06 PS=1.8e-06 $X=6060 $Y=1390 $dt=0
M7 9 15 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.95e-13 AS=1.659e-13 PD=2.23e-06 PS=1.21e-06 $X=7045 $Y=1390 $dt=0
M8 14 19 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=8695 $Y=1020 $dt=0
M9 13 9 14 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=9295 $Y=1020 $dt=0
M10 12 15 13 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=10185 $Y=1020 $dt=0
M11 8 11 12 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.55817e-13 AS=5.25e-14 PD=9.68244e-07 PS=6.7e-07 $X=10785 $Y=1020 $dt=0
M12 gnd3i! RN 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.60325e-13 AS=3.30183e-13 PD=1.475e-06 PS=2.05176e-06 $X=11755 $Y=660 $dt=0
M13 11 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=2.60325e-13 PD=2.74e-06 PS=1.475e-06 $X=12690 $Y=660 $dt=0
M14 Q 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=4.272e-13 PD=1.43e-06 PS=2.74e-06 $X=14280 $Y=660 $dt=0
M15 gnd3i! 13 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=15170 $Y=660 $dt=0
M16 Q 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=16060 $Y=660 $dt=0
M17 gnd3i! 13 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=2.403e-13 PD=2.74e-06 PS=1.43e-06 $X=16950 $Y=660 $dt=0
M18 vdd3i! 17 19 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.54046e-13 AS=6.768e-13 PD=2.58169e-06 PS=3.78e-06 $X=620 $Y=2410 $dt=1
M19 17 RN vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.136e-13 AS=2.31854e-13 PD=2.4e-06 PS=1.31831e-06 $X=1460 $Y=2670 $dt=1
M20 23 19 vdd3i! vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=5.1875e-13 PD=6.7e-07 PS=2.99e-06 $X=3080 $Y=3400 $dt=1
M21 17 15 23 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=1.21617e-13 AS=5.25e-14 PD=9.13043e-07 PS=6.7e-07 $X=3630 $Y=3400 $dt=1
M22 22 9 17 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=1.2e-13 AS=2.77983e-13 PD=1.21e-06 PS=2.08696e-06 $X=4470 $Y=2860 $dt=1
M23 vdd3i! D 22 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=5.00229e-13 AS=1.2e-13 PD=2.34286e-06 PS=1.21e-06 $X=5020 $Y=2860 $dt=1
M24 15 C vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=4.94875e-13 AS=3.75171e-13 PD=3.04e-06 PS=1.75714e-06 $X=6060 $Y=2860 $dt=1
M25 vdd3i! 15 9 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.92547e-13 AS=3.528e-13 PD=1.8586e-06 PS=2.42e-06 $X=7720 $Y=2670 $dt=1
M26 21 19 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=1.25e-13 AS=5.45203e-13 PD=1.25e-06 PS=2.5814e-06 $X=8740 $Y=2820 $dt=1
M27 13 15 21 vdd3i! pe3i L=3e-07 W=1e-06 AD=2.96338e-13 AS=1.25e-13 PD=2.19718e-06 PS=1.25e-06 $X=9290 $Y=2820 $dt=1
M28 20 9 13 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=1.24462e-13 PD=6.7e-07 PS=9.22817e-07 $X=10150 $Y=3235 $dt=1
M29 vdd3i! 11 20 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=2.90656e-13 AS=5.25e-14 PD=1.25671e-06 PS=6.7e-07 $X=10700 $Y=3235 $dt=1
M30 vdd3i! RN 13 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=4.98268e-13 AS=2.976e-13 PD=2.15435e-06 PS=2.4e-06 $X=11900 $Y=2410 $dt=1
M31 11 13 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=9.75775e-13 PD=3.78e-06 PS=4.21894e-06 $X=12740 $Y=2410 $dt=1
M32 Q 13 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=1.1618e-12 PD=1.95e-06 PS=4.88e-06 $X=14480 $Y=2410 $dt=1
M33 vdd3i! 13 Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=3.807e-13 PD=1.95e-06 PS=1.95e-06 $X=15320 $Y=2410 $dt=1
M34 Q 13 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=3.807e-13 PD=1.95e-06 PS=1.95e-06 $X=16160 $Y=2410 $dt=1
M35 vdd3i! 13 Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=3.807e-13 PD=3.78e-06 PS=1.95e-06 $X=17000 $Y=2410 $dt=1
.ends DFRRQJI3VX4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX0                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX0 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=4
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.923e-13 AS=2.016e-13 PD=2.005e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=3.923e-13 PD=1.8e-06 PS=2.005e-06 $X=1735 $Y=1130 $dt=0
M2 vdd3i! A 6 vdd3i! pe3i L=3e-07 W=9e-07 AD=5.7805e-13 AS=4.32e-13 PD=2.33911e-06 PS=2.76e-06 $X=620 $Y=2410 $dt=1
M3 Q 6 vdd3i! vdd3i! pe3i L=3e-07 W=1.12e-06 AD=5.376e-13 AS=7.1935e-13 PD=3.2e-06 PS=2.91089e-06 $X=1785 $Y=2410 $dt=1
.ends BUJI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AN21JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AN21JI3VX1 vdd3i! gnd3i! B A Q C
*.DEVICECLIMB
** N=9 EP=6 FDC=6
M0 8 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=6.47e-13 PD=1.14e-06 PS=3.58e-06 $X=690 $Y=660 $dt=0
M1 Q A 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.28413e-13 AS=1.1125e-13 PD=1.78572e-06 PS=1.14e-06 $X=1290 $Y=660 $dt=0
M2 gnd3i! C Q gnd3i! ne3i L=3.5e-07 W=6.65e-07 AD=6.369e-13 AS=2.45387e-13 PD=3.6e-06 PS=1.33428e-06 $X=2310 $Y=885 $dt=0
M3 vdd3i! B 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.371e-13 AS=6.768e-13 PD=2.03e-06 PS=3.78e-06 $X=620 $Y=2410 $dt=1
M4 9 A vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=4.371e-13 PD=1.95e-06 PS=2.03e-06 $X=1540 $Y=2410 $dt=1
M5 Q C 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.614e-13 AS=3.807e-13 PD=3.9e-06 PS=1.95e-06 $X=2380 $Y=2410 $dt=1
.ends AN21JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: EN3JI3VX1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt EN3JI3VX1 vdd3i! gnd3i! C B A Q
*.DEVICECLIMB
** N=16 EP=6 FDC=20
M0 13 C gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=2.016e-13 PD=9.6e-07 PS=1.8e-06 $X=620 $Y=1030 $dt=0
M1 gnd3i! B 13 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.97668e-13 AS=1.134e-13 PD=1.24213e-06 PS=9.6e-07 $X=1510 $Y=1030 $dt=0
M2 12 C gnd3i! gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=6.5e-14 AS=2.44732e-13 PD=7.7e-07 PS=1.53787e-06 $X=2730 $Y=930 $dt=0
M3 11 B 12 gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=1.404e-13 AS=6.5e-14 PD=1.06e-06 PS=7.7e-07 $X=3330 $Y=930 $dt=0
M4 gnd3i! 13 11 gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=5.308e-13 AS=1.404e-13 PD=3.32e-06 PS=1.06e-06 $X=4220 $Y=930 $dt=0
M5 9 11 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=5850 $Y=970 $dt=0
M6 gnd3i! A 9 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=6450 $Y=970 $dt=0
M7 8 A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=1.134e-13 PD=9.6e-07 PS=9.6e-07 $X=7340 $Y=970 $dt=0
M8 gnd3i! 11 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.965e-13 AS=1.134e-13 PD=3.17071e-06 PS=9.6e-07 $X=8230 $Y=970 $dt=0
M9 Q 10 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=2.0035e-13 PD=1.8e-06 PS=1.77071e-06 $X=9670 $Y=1130 $dt=0
M10 16 C vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.115e-13 AS=7.1585e-13 PD=1.71e-06 PS=3.85e-06 $X=645 $Y=2410 $dt=1
M11 13 B 16 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=5.5365e-13 AS=2.115e-13 PD=3.83e-06 PS=1.71e-06 $X=1245 $Y=2410 $dt=1
M12 vdd3i! C 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.23e-13 AS=5.8645e-13 PD=2.01e-06 PS=3.83e-06 $X=2675 $Y=2410 $dt=1
M13 14 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=4.23e-13 PD=2e-06 PS=2.01e-06 $X=3575 $Y=2410 $dt=1
M14 11 13 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.1205e-13 AS=4.1595e-13 PD=3.83e-06 PS=2e-06 $X=4465 $Y=2410 $dt=1
M15 10 11 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=9.1545e-13 PD=2e-06 PS=4.61e-06 $X=6095 $Y=2410 $dt=1
M16 vdd3i! A 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.956e-13 AS=4.1595e-13 PD=2.63e-06 PS=2e-06 $X=6985 $Y=2410 $dt=1
M17 15 A vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.115e-13 AS=6.956e-13 PD=1.71e-06 PS=2.63e-06 $X=8155 $Y=2410 $dt=1
M18 Q 11 15 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.66787e-13 AS=2.115e-13 PD=2.36668e-06 PS=1.71e-06 $X=8755 $Y=2410 $dt=1
M19 vdd3i! 10 Q vdd3i! pe3i L=3e-07 W=9.85e-07 AD=8.62325e-13 AS=3.26088e-13 PD=4.61e-06 PS=1.65332e-06 $X=9655 $Y=2410 $dt=1
.ends EN3JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA3I2JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA3I2JI3VX1 vdd3i! gnd3i! AN BN C Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 9 AN gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=4.00432e-13 PD=9.6e-07 PS=2.10243e-06 $X=540 $Y=1130 $dt=0
M1 gnd3i! BN 9 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=4.00432e-13 AS=1.134e-13 PD=2.10243e-06 PS=9.6e-07 $X=1430 $Y=1130 $dt=0
M2 8 C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=8.48535e-13 PD=1.14e-06 PS=4.45514e-06 $X=2290 $Y=660 $dt=0
M3 Q 9 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.806e-13 AS=1.1125e-13 PD=2.86e-06 PS=1.14e-06 $X=2890 $Y=660 $dt=0
M4 10 AN 9 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=4.08e-13 PD=1.1e-06 PS=2.66e-06 $X=620 $Y=2410 $dt=1
M5 vdd3i! BN 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=7.38476e-13 AS=1.0625e-13 PD=3.31526e-06 PS=1.1e-06 $X=1170 $Y=2410 $dt=1
M6 vdd3i! C Q vdd3i! pe3i L=3.00037e-07 W=1.00071e-06 AD=8.69412e-13 AS=2.376e-13 PD=3.90308e-06 PS=1.49071e-06 $X=2170 $Y=2410 $dt=1
M7 Q 9 vdd3i! vdd3i! pe3i L=3.00037e-07 W=1.00071e-06 AD=2.376e-13 AS=8.69412e-13 PD=1.49071e-06 PS=3.90308e-06 $X=3010 $Y=2410 $dt=1
.ends NA3I2JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA22JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA22JI3VX1 vdd3i! gnd3i! A B C Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 9 A 10 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=2.688e-13 PD=8.1e-07 PS=2.08e-06 $X=620 $Y=990 $dt=0
M1 gnd3i! B 9 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=3.3376e-13 AS=7e-14 PD=1.56028e-06 PS=8.1e-07 $X=1220 $Y=990 $dt=0
M2 8 C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=5.3044e-13 PD=1.14e-06 PS=2.47972e-06 $X=2350 $Y=660 $dt=0
M3 Q 10 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=1.1125e-13 PD=2.74e-06 PS=1.14e-06 $X=2950 $Y=660 $dt=0
M4 10 A vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=7.66562e-13 PD=1.24e-06 PS=3.33273e-06 $X=510 $Y=2410 $dt=1
M5 vdd3i! B 10 vdd3i! pe3i L=3e-07 W=7e-07 AD=7.66562e-13 AS=1.89e-13 PD=3.33273e-06 PS=1.24e-06 $X=1350 $Y=2410 $dt=1
M6 vdd3i! C Q vdd3i! pe3i L=3.00052e-07 W=9.98995e-07 AD=1.09399e-12 AS=2.255e-13 PD=4.75626e-06 PS=1.46899e-06 $X=2190 $Y=2410 $dt=1
M7 Q 10 vdd3i! vdd3i! pe3i L=3.00052e-07 W=9.98995e-07 AD=2.255e-13 AS=1.09399e-12 PD=1.46899e-06 PS=4.75626e-06 $X=3030 $Y=2410 $dt=1
.ends NA22JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AN22JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AN22JI3VX1 vdd3i! gnd3i! B A Q C D
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 10 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=6.098e-13 PD=1.14e-06 PS=3.52e-06 $X=660 $Y=660 $dt=0
M1 Q A 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=1.1125e-13 PD=1.43e-06 PS=1.14e-06 $X=1260 $Y=660 $dt=0
M2 9 C Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=2.403e-13 PD=1.14e-06 PS=1.43e-06 $X=2150 $Y=660 $dt=0
M3 gnd3i! D 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=8.082e-13 AS=1.1125e-13 PD=3.84e-06 PS=1.14e-06 $X=2750 $Y=660 $dt=0
M4 vdd3i! B 11 vdd3i! pe3i L=3.01094e-07 W=1.47213e-06 AD=4.29e-13 AS=6.0945e-13 PD=2.32213e-06 PS=3.77213e-06 $X=660 $Y=2410 $dt=1
M5 11 A vdd3i! vdd3i! pe3i L=3.01094e-07 W=1.47213e-06 AD=4.05825e-13 AS=4.29e-13 PD=2.06213e-06 PS=2.32213e-06 $X=1310 $Y=2410 $dt=1
M6 Q C 11 vdd3i! pe3i L=3.01094e-07 W=1.47213e-06 AD=2.9925e-13 AS=4.05825e-13 PD=1.92213e-06 PS=2.06213e-06 $X=2200 $Y=2410 $dt=1
M7 11 D Q vdd3i! pe3i L=3.01094e-07 W=1.47213e-06 AD=6.252e-13 AS=2.9925e-13 PD=3.77213e-06 PS=1.92213e-06 $X=3100 $Y=2410 $dt=1
.ends AN22JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DLY1JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DLY1JI3VX1 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=8 EP=4 FDC=8
M0 gnd3i! A 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.591e-13 AS=2.016e-13 PD=2.13e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 6 8 gnd3i! gnd3i! ne3i L=8e-07 W=4.2e-07 AD=2.415e-13 AS=3.591e-13 PD=1.99e-06 PS=2.13e-06 $X=1590 $Y=1400 $dt=0
M2 gnd3i! 6 7 gnd3i! ne3i L=1e-06 W=4.2e-07 AD=2.6662e-13 AS=2.016e-13 PD=1.28565e-06 PS=1.8e-06 $X=2860 $Y=660 $dt=0
M3 Q 7 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.3165e-13 AS=5.6498e-13 PD=2.75e-06 PS=2.72435e-06 $X=4625 $Y=660 $dt=0
M4 vdd3i! A 8 vdd3i! pe3i L=3e-07 W=6.7e-07 AD=4.61962e-13 AS=3.3835e-13 PD=2.62468e-06 PS=2.35e-06 $X=645 $Y=2680 $dt=1
M5 6 8 vdd3i! vdd3i! pe3i L=1e-06 W=4.2e-07 AD=2.00088e-13 AS=2.89588e-13 PD=1.76778e-06 PS=1.64532e-06 $X=1590 $Y=2680 $dt=1
M6 vdd3i! 6 7 vdd3i! pe3i L=7.5e-07 W=4.2e-07 AD=2.78313e-13 AS=2.00088e-13 PD=1.17049e-06 PS=1.76778e-06 $X=3110 $Y=3400 $dt=1
M7 Q 7 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.191e-13 AS=9.34337e-13 PD=3.84e-06 PS=3.92951e-06 $X=4650 $Y=2410 $dt=1
.ends DLY1JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ON21JI3VX4                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ON21JI3VX4 vdd3i! gnd3i! B A C Q
*.DEVICECLIMB
** N=11 EP=6 FDC=16
M0 gnd3i! B 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=4.272e-13 PD=1.43e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 10 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=1510 $Y=660 $dt=0
M2 9 C 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.868e-13 AS=2.403e-13 PD=2.70971e-06 PS=1.43e-06 $X=2400 $Y=660 $dt=0
M3 gnd3i! 9 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.35783e-13 AS=4.34e-13 PD=1.42065e-06 PS=2.92971e-06 $X=3930 $Y=660 $dt=0
M4 Q 8 gnd3i! gnd3i! ne3i L=3.49164e-07 W=8.96213e-07 AD=2.32912e-13 AS=2.37429e-13 PD=1.42121e-06 PS=1.43057e-06 $X=4820 $Y=660 $dt=0
M5 gnd3i! 8 Q gnd3i! ne3i L=3.49164e-07 W=8.96213e-07 AD=2.32912e-13 AS=2.32912e-13 PD=1.42121e-06 PS=1.42121e-06 $X=5680 $Y=660 $dt=0
M6 Q 8 gnd3i! gnd3i! ne3i L=3.49164e-07 W=8.96213e-07 AD=2.32912e-13 AS=2.32912e-13 PD=1.42121e-06 PS=1.42121e-06 $X=6570 $Y=660 $dt=0
M7 gnd3i! 8 Q gnd3i! ne3i L=3.49164e-07 W=8.96213e-07 AD=4.19812e-13 AS=2.32912e-13 PD=2.73121e-06 PS=1.42121e-06 $X=7430 $Y=660 $dt=0
M8 11 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=9.418e-13 PD=1.66e-06 PS=4.63e-06 $X=695 $Y=2410 $dt=1
M9 9 A 11 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.68825e-13 AS=1.7625e-13 PD=2.075e-06 PS=1.66e-06 $X=1245 $Y=2410 $dt=1
M10 vdd3i! C 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.285e-12 AS=4.68825e-13 PD=5.02e-06 PS=2.075e-06 $X=2210 $Y=2410 $dt=1
M11 vdd3i! 9 8 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=5.48179e-13 AS=6.768e-13 PD=2.4141e-06 PS=3.78e-06 $X=4020 $Y=2410 $dt=1
M12 Q 8 vdd3i! vdd3i! pe3i L=3.00021e-07 W=1.42657e-06 AD=3.433e-13 AS=5.54621e-13 PD=1.92657e-06 PS=2.44247e-06 $X=4960 $Y=2410 $dt=1
M13 vdd3i! 8 Q vdd3i! pe3i L=3.00021e-07 W=1.42657e-06 AD=4.866e-13 AS=3.433e-13 PD=2.35657e-06 PS=1.92657e-06 $X=5800 $Y=2410 $dt=1
M14 Q 8 vdd3i! vdd3i! pe3i L=3.00021e-07 W=1.42657e-06 AD=3.433e-13 AS=4.866e-13 PD=1.92657e-06 PS=2.35657e-06 $X=6640 $Y=2410 $dt=1
M15 vdd3i! 8 Q vdd3i! pe3i L=3.00021e-07 W=1.42657e-06 AD=8.562e-13 AS=3.433e-13 PD=4.53657e-06 PS=1.92657e-06 $X=7480 $Y=2410 $dt=1
.ends ON21JI3VX4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INJI3VX6                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INJI3VX6 vdd3i! gnd3i! Q A
*.DEVICECLIMB
** N=5 EP=4 FDC=10
M0 gnd3i! A Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=4.272e-13 PD=1.86e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=1590 $Y=660 $dt=0
M2 gnd3i! A Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.114e-13 AS=2.403e-13 PD=1.96e-06 PS=1.43e-06 $X=2480 $Y=660 $dt=0
M3 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=4.114e-13 PD=2.74e-06 PS=1.96e-06 $X=3550 $Y=660 $dt=0
M4 Q A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=5.79287e-13 PD=1.86506e-06 PS=3.69506e-06 $X=475 $Y=2410 $dt=1
M5 vdd3i! A Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1315 $Y=2410 $dt=1
M6 Q A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1865 $Y=2410 $dt=1
M7 vdd3i! A Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=2705 $Y=2410 $dt=1
M8 Q A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=3255 $Y=2410 $dt=1
M9 vdd3i! A Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=1.01149e-12 AS=2.54913e-13 PD=4.73506e-06 PS=1.86506e-06 $X=4095 $Y=2410 $dt=1
.ends INJI3VX6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA3I1JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA3I1JI3VX1 vdd3i! gnd3i! AN Q B C
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 gnd3i! AN 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.40779e-13 AS=2.016e-13 PD=1.24397e-06 PS=1.8e-06 $X=620 $Y=660 $dt=0
M1 9 10 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.26825e-13 AS=5.10221e-13 PD=1.175e-06 PS=2.63603e-06 $X=1670 $Y=660 $dt=0
M2 8 B 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.31275e-13 AS=1.26825e-13 PD=1.185e-06 PS=1.175e-06 $X=2305 $Y=660 $dt=0
M3 Q C 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=1.31275e-13 PD=2.74e-06 PS=1.185e-06 $X=2950 $Y=660 $dt=0
M4 vdd3i! AN 10 vdd3i! pe3i L=3e-07 W=7e-07 AD=4.82246e-13 AS=3.36e-13 PD=2.26063e-06 PS=2.36e-06 $X=620 $Y=2410 $dt=1
M5 vdd3i! 10 Q vdd3i! pe3i L=3.00059e-07 W=1.00314e-06 AD=6.91085e-13 AS=2.195e-13 PD=3.2396e-06 PS=1.46314e-06 $X=1430 $Y=2410 $dt=1
M6 Q B vdd3i! vdd3i! pe3i L=3.00059e-07 W=1.00314e-06 AD=2.195e-13 AS=6.91085e-13 PD=1.46314e-06 PS=3.2396e-06 $X=2270 $Y=2410 $dt=1
M7 Q C vdd3i! vdd3i! pe3i L=3.00059e-07 W=1.00314e-06 AD=4.232e-13 AS=6.91085e-13 PD=2.85314e-06 PS=3.2396e-06 $X=3000 $Y=2410 $dt=1
.ends NA3I1JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX8                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX8 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=19
M0 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=6.098e-13 PD=1.43e-06 PS=3.52e-06 $X=660 $Y=660 $dt=0
M1 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.804e-13 AS=2.403e-13 PD=1.91e-06 PS=1.43e-06 $X=1550 $Y=660 $dt=0
M2 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.804e-13 PD=1.43e-06 PS=1.91e-06 $X=2570 $Y=660 $dt=0
M3 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=3460 $Y=660 $dt=0
M4 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=4430 $Y=660 $dt=0
M5 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=5320 $Y=660 $dt=0
M6 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=6290 $Y=660 $dt=0
M7 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=8.702e-13 AS=2.403e-13 PD=3.94e-06 PS=1.43e-06 $X=7180 $Y=660 $dt=0
M8 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=5.51013e-13 PD=1.86506e-06 PS=3.69506e-06 $X=620 $Y=2410 $dt=1
M9 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.61963e-13 AS=2.83187e-13 PD=1.87506e-06 PS=1.86506e-06 $X=1170 $Y=2410 $dt=1
M10 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.61963e-13 PD=1.86506e-06 PS=1.87506e-06 $X=2020 $Y=2410 $dt=1
M11 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.61963e-13 AS=2.83187e-13 PD=1.87506e-06 PS=1.86506e-06 $X=2570 $Y=2410 $dt=1
M12 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.61963e-13 PD=1.86506e-06 PS=1.87506e-06 $X=3420 $Y=2410 $dt=1
M13 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.61963e-13 AS=2.83187e-13 PD=1.87506e-06 PS=1.86506e-06 $X=3970 $Y=2410 $dt=1
M14 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.61963e-13 PD=1.86506e-06 PS=1.87506e-06 $X=4820 $Y=2410 $dt=1
M15 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.61963e-13 AS=2.83187e-13 PD=1.87506e-06 PS=1.86506e-06 $X=5370 $Y=2410 $dt=1
M16 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.61963e-13 PD=1.86506e-06 PS=1.87506e-06 $X=6220 $Y=2410 $dt=1
M17 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.61963e-13 AS=2.83187e-13 PD=1.87506e-06 PS=1.86506e-06 $X=6770 $Y=2410 $dt=1
M18 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=5.79287e-13 AS=2.61963e-13 PD=3.69506e-06 PS=1.87506e-06 $X=7620 $Y=2410 $dt=1
.ends BUJI3VX8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DFRRQJI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DFRRQJI3VX1 vdd3i! gnd3i! RN D C Q
*.DEVICECLIMB
** N=23 EP=6 FDC=30
M0 gnd3i! 17 19 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.39017e-13 AS=2.016e-13 PD=9.16947e-07 PS=1.8e-06 $X=620 $Y=660 $dt=0
M1 10 RN gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.28952e-13 AS=2.94583e-13 PD=2.36956e-06 PS=1.94305e-06 $X=1510 $Y=660 $dt=0
M2 18 19 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.55236e-13 PD=6.7e-07 PS=1.11822e-06 $X=2340 $Y=1390 $dt=0
M3 17 9 18 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=2940 $Y=1390 $dt=0
M4 16 15 17 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=3830 $Y=1390 $dt=0
M5 10 D 16 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.835e-13 AS=5.25e-14 PD=2.19e-06 PS=6.7e-07 $X=4430 $Y=1390 $dt=0
M6 gnd3i! C 15 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.659e-13 AS=2.016e-13 PD=1.21e-06 PS=1.8e-06 $X=6060 $Y=1390 $dt=0
M7 9 15 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.95e-13 AS=1.659e-13 PD=2.23e-06 PS=1.21e-06 $X=7045 $Y=1390 $dt=0
M8 14 19 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=8695 $Y=1020 $dt=0
M9 13 9 14 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=9295 $Y=1020 $dt=0
M10 12 15 13 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=10185 $Y=1020 $dt=0
M11 8 11 12 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.55817e-13 AS=5.25e-14 PD=9.68244e-07 PS=6.7e-07 $X=10785 $Y=1020 $dt=0
M12 gnd3i! RN 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=6.52289e-13 AS=3.30183e-13 PD=3.3375e-06 PS=2.05176e-06 $X=11755 $Y=660 $dt=0
M13 11 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=3.07822e-13 PD=1.8e-06 PS=1.575e-06 $X=12560 $Y=1130 $dt=0
M14 Q 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=6.52289e-13 PD=2.74e-06 PS=3.3375e-06 $X=14150 $Y=660 $dt=0
M15 vdd3i! 17 19 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=1.944e-13 AS=3.456e-13 PD=1.26e-06 PS=2.4e-06 $X=620 $Y=2670 $dt=1
M16 17 RN vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.136e-13 AS=1.944e-13 PD=2.4e-06 PS=1.26e-06 $X=1460 $Y=2670 $dt=1
M17 23 19 vdd3i! vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=5.1875e-13 PD=6.7e-07 PS=2.99e-06 $X=3080 $Y=3400 $dt=1
M18 17 15 23 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=1.21617e-13 AS=5.25e-14 PD=9.13043e-07 PS=6.7e-07 $X=3630 $Y=3400 $dt=1
M19 22 9 17 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=1.2e-13 AS=2.77983e-13 PD=1.21e-06 PS=2.08696e-06 $X=4470 $Y=2860 $dt=1
M20 vdd3i! D 22 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=5.00229e-13 AS=1.2e-13 PD=2.34286e-06 PS=1.21e-06 $X=5020 $Y=2860 $dt=1
M21 15 C vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=4.94875e-13 AS=3.75171e-13 PD=3.04e-06 PS=1.75714e-06 $X=6060 $Y=2860 $dt=1
M22 vdd3i! 15 9 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.92547e-13 AS=3.528e-13 PD=1.8586e-06 PS=2.42e-06 $X=7720 $Y=2670 $dt=1
M23 21 19 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=1.25e-13 AS=5.45203e-13 PD=1.25e-06 PS=2.5814e-06 $X=8740 $Y=2820 $dt=1
M24 13 15 21 vdd3i! pe3i L=3e-07 W=1e-06 AD=2.96338e-13 AS=1.25e-13 PD=2.19718e-06 PS=1.25e-06 $X=9290 $Y=2820 $dt=1
M25 20 9 13 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=1.24462e-13 PD=6.7e-07 PS=9.22817e-07 $X=10150 $Y=3235 $dt=1
M26 vdd3i! 11 20 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=4.10996e-13 AS=5.25e-14 PD=1.64789e-06 PS=6.7e-07 $X=10700 $Y=3235 $dt=1
M27 vdd3i! RN 13 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=7.04565e-13 AS=2.976e-13 PD=2.82495e-06 PS=2.4e-06 $X=11900 $Y=2410 $dt=1
M28 11 13 vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.456e-13 AS=7.04565e-13 PD=2.4e-06 PS=2.82495e-06 $X=12740 $Y=2410 $dt=1
M29 Q 13 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=1.37977e-12 PD=3.78e-06 PS=5.5322e-06 $X=14200 $Y=2410 $dt=1
.ends DFRRQJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ON211JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ON211JI3VX1 vdd3i! gnd3i! B Q A C D
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 Q B 10 gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.27987e-13 AS=4.20337e-13 PD=1.41536e-06 PS=2.75536e-06 $X=620 $Y=660 $dt=0
M1 10 A Q gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.30287e-13 AS=2.27987e-13 PD=1.43036e-06 PS=1.41536e-06 $X=1460 $Y=660 $dt=0
M2 9 C 10 gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=1.21188e-13 AS=2.30287e-13 PD=1.17536e-06 PS=1.43036e-06 $X=2350 $Y=660 $dt=0
M3 gnd3i! D 9 gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=4.20337e-13 AS=1.21188e-13 PD=2.75536e-06 PS=1.17536e-06 $X=2950 $Y=660 $dt=0
M4 11 B vdd3i! vdd3i! pe3i L=3e-07 W=1.38e-06 AD=1.725e-13 AS=9.388e-13 PD=1.63e-06 PS=4.63e-06 $X=695 $Y=2410 $dt=1
M5 Q A 11 vdd3i! pe3i L=3e-07 W=1.38e-06 AD=4.69617e-13 AS=1.725e-13 PD=2.38255e-06 PS=1.63e-06 $X=1245 $Y=2410 $dt=1
M6 vdd3i! C Q vdd3i! pe3i L=3.00049e-07 W=9.66924e-07 AD=4.25413e-13 AS=3.29046e-13 PD=2.34192e-06 PS=1.66938e-06 $X=2210 $Y=2410 $dt=1
M7 Q D vdd3i! vdd3i! pe3i L=3.00049e-07 W=9.66924e-07 AD=4.20162e-13 AS=4.25413e-13 PD=2.80192e-06 PS=2.34192e-06 $X=3000 $Y=2410 $dt=1
.ends ON211JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ON22JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ON22JI3VX1 vdd3i! gnd3i! D C Q A B
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 gnd3i! D 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=4.272e-13 PD=1.86e-06 PS=2.74e-06 $X=720 $Y=660 $dt=0
M1 9 C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=1690 $Y=660 $dt=0
M2 Q A 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=2580 $Y=660 $dt=0
M3 9 B Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.666e-13 AS=2.403e-13 PD=2.84e-06 PS=1.43e-06 $X=3470 $Y=660 $dt=0
M4 11 D vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=8.802e-13 PD=1.66e-06 PS=4.56e-06 $X=1120 $Y=2410 $dt=1
M5 Q C 11 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=1.7625e-13 PD=1.95e-06 PS=1.66e-06 $X=1670 $Y=2410 $dt=1
M6 10 A Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=3.807e-13 PD=1.66e-06 PS=1.95e-06 $X=2510 $Y=2410 $dt=1
M7 vdd3i! B 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=8.802e-13 AS=1.7625e-13 PD=4.56e-06 PS=1.66e-06 $X=3060 $Y=2410 $dt=1
.ends ON22JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DFRRQJI3VX2                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DFRRQJI3VX2 vdd3i! gnd3i! RN D C Q
*.DEVICECLIMB
** N=23 EP=6 FDC=32
M0 gnd3i! 17 19 gnd3i! ne3i L=3.5e-07 W=6.6e-07 AD=1.94849e-13 AS=3.168e-13 PD=1.21781e-06 PS=2.28e-06 $X=620 $Y=660 $dt=0
M1 10 RN gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.28952e-13 AS=2.62751e-13 PD=2.36956e-06 PS=1.64219e-06 $X=1510 $Y=660 $dt=0
M2 18 19 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.55236e-13 PD=6.7e-07 PS=1.11822e-06 $X=2340 $Y=1390 $dt=0
M3 17 9 18 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=2940 $Y=1390 $dt=0
M4 16 15 17 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=3830 $Y=1390 $dt=0
M5 10 D 16 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.835e-13 AS=5.25e-14 PD=2.19e-06 PS=6.7e-07 $X=4430 $Y=1390 $dt=0
M6 gnd3i! C 15 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.659e-13 AS=2.016e-13 PD=1.21e-06 PS=1.8e-06 $X=6060 $Y=1390 $dt=0
M7 9 15 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.95e-13 AS=1.659e-13 PD=2.23e-06 PS=1.21e-06 $X=7045 $Y=1390 $dt=0
M8 14 19 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=8695 $Y=1020 $dt=0
M9 13 9 14 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=9295 $Y=1020 $dt=0
M10 12 15 13 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=10185 $Y=1020 $dt=0
M11 8 11 12 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.55817e-13 AS=5.25e-14 PD=9.68244e-07 PS=6.7e-07 $X=10785 $Y=1020 $dt=0
M12 gnd3i! RN 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=5.94987e-13 AS=3.30183e-13 PD=3.35209e-06 PS=2.05176e-06 $X=11755 $Y=660 $dt=0
M13 11 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=6.6e-07 AD=3.168e-13 AS=4.41226e-13 PD=2.28e-06 PS=2.48582e-06 $X=12750 $Y=890 $dt=0
M14 Q 13 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=5.94987e-13 PD=1.43e-06 PS=3.35209e-06 $X=14380 $Y=660 $dt=0
M15 gnd3i! 13 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=2.403e-13 PD=2.74e-06 PS=1.43e-06 $X=15270 $Y=660 $dt=0
M16 vdd3i! 17 19 vdd3i! pe3i L=3e-07 W=1e-06 AD=2.97674e-13 AS=4.8e-13 PD=1.7907e-06 PS=2.96e-06 $X=620 $Y=2670 $dt=1
M17 17 RN vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.136e-13 AS=2.14326e-13 PD=2.4e-06 PS=1.2893e-06 $X=1460 $Y=2670 $dt=1
M18 23 19 vdd3i! vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=5.1875e-13 PD=6.7e-07 PS=2.99e-06 $X=3080 $Y=3400 $dt=1
M19 17 15 23 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=1.21617e-13 AS=5.25e-14 PD=9.13043e-07 PS=6.7e-07 $X=3630 $Y=3400 $dt=1
M20 22 9 17 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=1.2e-13 AS=2.77983e-13 PD=1.21e-06 PS=2.08696e-06 $X=4470 $Y=2860 $dt=1
M21 vdd3i! D 22 vdd3i! pe3i L=3e-07 W=9.6e-07 AD=5.00229e-13 AS=1.2e-13 PD=2.34286e-06 PS=1.21e-06 $X=5020 $Y=2860 $dt=1
M22 15 C vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=4.56625e-13 AS=3.75171e-13 PD=2.86e-06 PS=1.75714e-06 $X=6060 $Y=2860 $dt=1
M23 vdd3i! 15 9 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.92547e-13 AS=3.528e-13 PD=1.8586e-06 PS=2.42e-06 $X=7720 $Y=2670 $dt=1
M24 21 19 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=1.25e-13 AS=5.45203e-13 PD=1.25e-06 PS=2.5814e-06 $X=8740 $Y=2820 $dt=1
M25 13 15 21 vdd3i! pe3i L=3e-07 W=1e-06 AD=2.96338e-13 AS=1.25e-13 PD=2.19718e-06 PS=1.25e-06 $X=9290 $Y=2820 $dt=1
M26 20 9 13 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=1.24462e-13 PD=6.7e-07 PS=9.22817e-07 $X=10150 $Y=3235 $dt=1
M27 vdd3i! 11 20 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=3.93439e-13 AS=5.25e-14 PD=1.64096e-06 PS=6.7e-07 $X=10700 $Y=3235 $dt=1
M28 vdd3i! RN 13 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=6.74468e-13 AS=2.976e-13 PD=2.81307e-06 PS=2.4e-06 $X=11900 $Y=2410 $dt=1
M29 11 13 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=4.8e-13 AS=9.36761e-13 PD=2.96e-06 PS=3.90704e-06 $X=12740 $Y=2410 $dt=1
M30 Q 13 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=1.32083e-12 PD=1.95e-06 PS=5.50893e-06 $X=14440 $Y=2410 $dt=1
M31 vdd3i! 13 Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=8.802e-13 AS=3.807e-13 PD=4.56e-06 PS=1.95e-06 $X=15280 $Y=2410 $dt=1
.ends DFRRQJI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: EO3JI3VX1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt EO3JI3VX1 vdd3i! gnd3i! C B A Q
*.DEVICECLIMB
** N=16 EP=6 FDC=20
M0 12 C gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.628e-13 PD=9.6e-07 PS=3.52e-06 $X=660 $Y=1130 $dt=0
M1 gnd3i! B 12 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.30196e-13 AS=1.134e-13 PD=1.36723e-06 PS=9.6e-07 $X=1550 $Y=1130 $dt=0
M2 11 C gnd3i! gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=6.5e-14 AS=2.85004e-13 PD=7.7e-07 PS=1.69277e-06 $X=2910 $Y=1030 $dt=0
M3 10 B 11 gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=1.404e-13 AS=6.5e-14 PD=1.06e-06 PS=7.7e-07 $X=3510 $Y=1030 $dt=0
M4 gnd3i! 12 10 gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=8.05779e-13 AS=1.404e-13 PD=2.83787e-06 PS=1.06e-06 $X=4400 $Y=1030 $dt=0
M5 9 10 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=6.50821e-13 PD=9.6e-07 PS=2.29213e-06 $X=6075 $Y=1130 $dt=0
M6 gnd3i! A 9 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.90537e-13 AS=1.134e-13 PD=1.53255e-06 PS=9.6e-07 $X=6965 $Y=1130 $dt=0
M7 8 A gnd3i! gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=6.5e-14 AS=3.59713e-13 PD=7.7e-07 PS=1.89745e-06 $X=8140 $Y=1030 $dt=0
M8 Q 10 8 gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=1.404e-13 AS=6.5e-14 PD=1.06e-06 PS=7.7e-07 $X=8740 $Y=1030 $dt=0
M9 gnd3i! 9 Q gnd3i! ne3i L=3.5e-07 W=5.2e-07 AD=5.728e-13 AS=1.404e-13 PD=3.52e-06 PS=1.06e-06 $X=9630 $Y=1030 $dt=0
M10 16 C vdd3i! vdd3i! pe3i L=3e-07 W=1.3e-06 AD=1.95e-13 AS=6.603e-13 PD=1.6e-06 PS=3.63e-06 $X=645 $Y=2520 $dt=1
M11 12 B 16 vdd3i! pe3i L=3e-07 W=1.3e-06 AD=5.157e-13 AS=1.95e-13 PD=3.61e-06 PS=1.6e-06 $X=1245 $Y=2520 $dt=1
M12 vdd3i! C 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=5.8645e-13 PD=2e-06 PS=3.83e-06 $X=2675 $Y=2410 $dt=1
M13 14 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=4.1595e-13 PD=2e-06 PS=2e-06 $X=3565 $Y=2410 $dt=1
M14 10 12 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=5.6965e-13 AS=4.1595e-13 PD=3.83e-06 PS=2e-06 $X=4455 $Y=2410 $dt=1
M15 15 10 vdd3i! vdd3i! pe3i L=3e-07 W=1.3e-06 AD=1.95e-13 AS=5.301e-13 PD=1.6e-06 PS=3.61e-06 $X=5885 $Y=2410 $dt=1
M16 9 A 15 vdd3i! pe3i L=3e-07 W=1.3e-06 AD=5.157e-13 AS=1.95e-13 PD=3.61e-06 PS=1.6e-06 $X=6485 $Y=2410 $dt=1
M17 vdd3i! A 13 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=5.8645e-13 PD=2e-06 PS=3.83e-06 $X=7915 $Y=2410 $dt=1
M18 13 10 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=4.1595e-13 PD=2e-06 PS=2e-06 $X=8805 $Y=2410 $dt=1
M19 Q 9 13 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.1205e-13 AS=4.1595e-13 PD=3.83e-06 PS=2e-06 $X=9695 $Y=2410 $dt=1
.ends EO3JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO2JI3VX0 vdd3i! gnd3i! B Q A
*.DEVICECLIMB
** N=7 EP=5 FDC=4
M0 Q B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=7.244e-13 PD=9.6e-07 PS=4.14e-06 $X=500 $Y=1130 $dt=0
M1 gnd3i! A Q gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=7.244e-13 AS=1.134e-13 PD=4.14e-06 PS=9.6e-07 $X=1390 $Y=1130 $dt=0
M2 7 B vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=9.298e-13 PD=1.1e-06 PS=4.68e-06 $X=720 $Y=2410 $dt=1
M3 Q A 7 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.08e-13 AS=1.0625e-13 PD=2.66e-06 PS=1.1e-06 $X=1270 $Y=2410 $dt=1
.ends NO2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ON21JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ON21JI3VX1 vdd3i! gnd3i! B A Q C
*.DEVICECLIMB
** N=9 EP=6 FDC=6
M0 gnd3i! B 8 gnd3i! ne3i L=3.4958e-07 W=8.92071e-07 AD=2.40125e-13 AS=4.24712e-13 PD=1.43207e-06 PS=2.73707e-06 $X=615 $Y=660 $dt=0
M1 8 A gnd3i! gnd3i! ne3i L=3.4958e-07 W=8.92071e-07 AD=2.37987e-13 AS=2.40125e-13 PD=1.42707e-06 PS=1.43207e-06 $X=1505 $Y=660 $dt=0
M2 Q C 8 gnd3i! ne3i L=3.4958e-07 W=8.92071e-07 AD=4.24712e-13 AS=2.37987e-13 PD=2.73707e-06 PS=1.42707e-06 $X=2395 $Y=660 $dt=0
M3 9 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=9.418e-13 PD=1.66e-06 PS=4.63e-06 $X=695 $Y=2410 $dt=1
M4 Q A 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.75706e-13 AS=1.7625e-13 PD=2.44322e-06 PS=1.66e-06 $X=1245 $Y=2410 $dt=1
M5 vdd3i! C Q vdd3i! pe3i L=3e-07 W=9.85e-07 AD=1.1721e-12 AS=3.32319e-13 PD=4.94e-06 PS=1.70678e-06 $X=2210 $Y=2410 $dt=1
.ends ON21JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OR4JI3VX1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OR4JI3VX1 vdd3i! gnd3i! C D Q B A
*.DEVICECLIMB
** N=13 EP=7 FDC=12
M0 11 C gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=4.12474e-13 PD=9.6e-07 PS=2.12185e-06 $X=510 $Y=1130 $dt=0
M1 gnd3i! D 11 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=4.12474e-13 AS=1.134e-13 PD=2.12185e-06 PS=9.6e-07 $X=1400 $Y=1130 $dt=0
M2 10 11 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=8.74052e-13 PD=1.14e-06 PS=4.4963e-06 $X=2330 $Y=660 $dt=0
M3 Q 9 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.56e-13 AS=1.1125e-13 PD=2.64627e-06 PS=1.14e-06 $X=2930 $Y=660 $dt=0
M4 9 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=7.908e-13 PD=9.6e-07 PS=4.27314e-06 $X=4410 $Y=1130 $dt=0
M5 gnd3i! A 9 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=7.908e-13 AS=1.134e-13 PD=4.27314e-06 PS=9.6e-07 $X=5300 $Y=1130 $dt=0
M6 13 C 11 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=4.08e-13 PD=1.1e-06 PS=2.66e-06 $X=620 $Y=2410 $dt=1
M7 vdd3i! D 13 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=6.21177e-13 AS=1.0625e-13 PD=2.08363e-06 PS=1.1e-06 $X=1170 $Y=2410 $dt=1
M8 Q 11 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=1.03042e-12 PD=1.95e-06 PS=3.45637e-06 $X=2480 $Y=2410 $dt=1
M9 vdd3i! 9 Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.09631e-12 AS=3.807e-13 PD=3.53124e-06 PS=1.95e-06 $X=3320 $Y=2410 $dt=1
M10 12 B vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=6.60894e-13 PD=1.1e-06 PS=2.12876e-06 $X=4690 $Y=2410 $dt=1
M11 9 A 12 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.08e-13 AS=1.0625e-13 PD=2.66e-06 PS=1.1e-06 $X=5240 $Y=2410 $dt=1
.ends OR4JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX16                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX16 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=39
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=4.272e-13 PD=1.43e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=1510 $Y=660 $dt=0
M2 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=2400 $Y=660 $dt=0
M3 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=3290 $Y=660 $dt=0
M4 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=2.403e-13 PD=1.43e-06 PS=1.43e-06 $X=4180 $Y=660 $dt=0
M5 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.4475e-13 AS=2.403e-13 PD=1.44e-06 PS=1.43e-06 $X=5070 $Y=660 $dt=0
M6 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.63267e-13 AS=2.4475e-13 PD=1.95905e-06 PS=1.44e-06 $X=5970 $Y=660 $dt=0
M7 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.26533e-13 PD=1.34e-06 PS=1.76095e-06 $X=6940 $Y=750 $dt=0
M8 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=7830 $Y=750 $dt=0
M9 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=8800 $Y=750 $dt=0
M10 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=9690 $Y=750 $dt=0
M11 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=10660 $Y=750 $dt=0
M12 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=11550 $Y=750 $dt=0
M13 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=12520 $Y=750 $dt=0
M14 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=13410 $Y=750 $dt=0
M15 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=14380 $Y=750 $dt=0
M16 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.84e-13 AS=2.16e-13 PD=2.56e-06 PS=1.34e-06 $X=15270 $Y=750 $dt=0
M17 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=5.79287e-13 PD=1.86506e-06 PS=3.69506e-06 $X=475 $Y=2410 $dt=1
M18 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1315 $Y=2410 $dt=1
M19 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1865 $Y=2410 $dt=1
M20 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=2705 $Y=2410 $dt=1
M21 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=3255 $Y=2410 $dt=1
M22 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=4095 $Y=2410 $dt=1
M23 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=4645 $Y=2410 $dt=1
M24 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=5485 $Y=2410 $dt=1
M25 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=6035 $Y=2410 $dt=1
M26 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=6875 $Y=2410 $dt=1
M27 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=7425 $Y=2410 $dt=1
M28 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=8265 $Y=2410 $dt=1
M29 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=8815 $Y=2410 $dt=1
M30 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=9655 $Y=2410 $dt=1
M31 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=10205 $Y=2410 $dt=1
M32 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=11045 $Y=2410 $dt=1
M33 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=11595 $Y=2410 $dt=1
M34 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=12435 $Y=2410 $dt=1
M35 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=12985 $Y=2410 $dt=1
M36 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=13825 $Y=2410 $dt=1
M37 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=14375 $Y=2410 $dt=1
M38 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=1.15229e-12 AS=2.54913e-13 PD=4.89506e-06 PS=1.86506e-06 $X=15215 $Y=2410 $dt=1
.ends BUJI3VX16

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX6                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX6 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=14
M0 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=6.008e-13 PD=1.34e-06 PS=3.52e-06 $X=660 $Y=750 $dt=0
M1 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=5.84805e-13 AS=2.16e-13 PD=2.17751e-06 PS=1.34e-06 $X=1550 $Y=750 $dt=0
M2 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=6.50595e-13 PD=1.43e-06 PS=2.42249e-06 $X=2960 $Y=660 $dt=0
M3 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=3850 $Y=660 $dt=0
M4 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=4820 $Y=660 $dt=0
M5 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=6.098e-13 AS=2.403e-13 PD=3.52e-06 PS=1.43e-06 $X=5710 $Y=660 $dt=0
M6 6 A vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=6.3285e-13 PD=1.87971e-06 PS=3.75971e-06 $X=525 $Y=2410 $dt=1
M7 vdd3i! A 6 vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=3.7905e-13 AS=2.751e-13 PD=1.98971e-06 PS=1.87971e-06 $X=1365 $Y=2410 $dt=1
M8 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=3.7905e-13 PD=1.87971e-06 PS=1.98971e-06 $X=2075 $Y=2410 $dt=1
M9 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=3.3675e-13 AS=2.751e-13 PD=1.92971e-06 PS=1.87971e-06 $X=2915 $Y=2410 $dt=1
M10 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=3.3675e-13 PD=1.87971e-06 PS=1.92971e-06 $X=3565 $Y=2410 $dt=1
M11 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=3.3675e-13 AS=2.751e-13 PD=1.92971e-06 PS=1.87971e-06 $X=4405 $Y=2410 $dt=1
M12 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=3.3675e-13 PD=1.87971e-06 PS=1.92971e-06 $X=5055 $Y=2410 $dt=1
M13 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=6.3285e-13 AS=2.751e-13 PD=3.75971e-06 PS=1.87971e-06 $X=5895 $Y=2410 $dt=1
.ends BUJI3VX6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ON31JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ON31JI3VX1 vdd3i! gnd3i! A B C Q D
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 9 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=6.098e-13 PD=1.43e-06 PS=3.52e-06 $X=660 $Y=660 $dt=0
M1 gnd3i! B 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=1550 $Y=660 $dt=0
M2 9 C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=2520 $Y=660 $dt=0
M3 Q D 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=2.403e-13 PD=2.74e-06 PS=1.43e-06 $X=3410 $Y=660 $dt=0
M4 11 A vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=9.066e-13 PD=1.72e-06 PS=4.59e-06 $X=1145 $Y=2410 $dt=1
M5 10 B 11 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=2.1855e-13 PD=1.72e-06 PS=1.72e-06 $X=1755 $Y=2410 $dt=1
M6 Q C 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=5.30442e-13 AS=2.1855e-13 PD=2.60067e-06 PS=1.72e-06 $X=2365 $Y=2410 $dt=1
M7 vdd3i! D Q vdd3i! pe3i L=3e-07 W=8.4e-07 AD=1.1576e-12 AS=3.16008e-13 PD=4.94e-06 PS=1.54933e-06 $X=3330 $Y=2410 $dt=1
.ends ON31JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DLY4JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DLY4JI3VX1 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=12 EP=4 FDC=12
M0 gnd3i! A 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.323e-13 AS=2.016e-13 PD=1.05e-06 PS=1.8e-06 $X=620 $Y=660 $dt=0
M1 8 10 gnd3i! gnd3i! ne3i L=1.8e-06 W=4.2e-07 AD=1.736e-13 AS=1.323e-13 PD=1.58e-06 PS=1.05e-06 $X=1600 $Y=660 $dt=0
M2 8 10 9 gnd3i! ne3i L=1.8e-06 W=4.2e-07 AD=1.736e-13 AS=2.00088e-13 PD=1.58e-06 PS=1.76778e-06 $X=1600 $Y=1360 $dt=0
M3 gnd3i! 9 7 gnd3i! ne3i L=1.1e-06 W=4.2e-07 AD=4.30324e-13 AS=2.16e-13 PD=1.75053e-06 PS=1.66e-06 $X=4630 $Y=660 $dt=0
M4 6 9 7 gnd3i! ne3i L=1.1e-06 W=4.2e-07 AD=2.00088e-13 AS=2.16e-13 PD=1.76778e-06 PS=1.66e-06 $X=4630 $Y=1400 $dt=0
M5 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.4055e-13 AS=9.11876e-13 PD=2.77e-06 PS=3.70947e-06 $X=7220 $Y=660 $dt=0
M6 vdd3i! A 10 vdd3i! pe3i L=3e-07 W=7e-07 AD=5.26875e-13 AS=3.535e-13 PD=3.30625e-06 PS=2.41e-06 $X=645 $Y=2680 $dt=1
M7 12 10 9 vdd3i! pe3i L=1.2e-06 W=4.2e-07 AD=1.674e-13 AS=2.016e-13 PD=1.56e-06 PS=1.8e-06 $X=2100 $Y=2680 $dt=1
M8 12 10 vdd3i! vdd3i! pe3i L=1.2e-06 W=4.2e-07 AD=1.674e-13 AS=3.16125e-13 PD=1.56e-06 PS=1.98375e-06 $X=2100 $Y=3400 $dt=1
M9 6 9 11 vdd3i! pe3i L=1.9e-06 W=4.2e-07 AD=2.016e-13 AS=1.674e-13 PD=1.8e-06 PS=1.56e-06 $X=4220 $Y=2680 $dt=1
M10 vdd3i! 9 11 vdd3i! pe3i L=1.9e-06 W=4.2e-07 AD=2.6367e-13 AS=1.674e-13 PD=1.32426e-06 PS=1.56e-06 $X=4220 $Y=3400 $dt=1
M11 Q 6 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.332e-13 AS=8.8518e-13 PD=3.86e-06 PS=4.44574e-06 $X=7245 $Y=2410 $dt=1
.ends DLY4JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO2I1JI3VX2                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO2I1JI3VX2 vdd3i! gnd3i! AN Q B
*.DEVICECLIMB
** N=9 EP=5 FDC=10
M0 gnd3i! AN 7 gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.3695e-13 AS=4.15012e-13 PD=1.44536e-06 PS=2.72536e-06 $X=595 $Y=660 $dt=0
M1 Q 7 gnd3i! gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.28113e-13 AS=2.3695e-13 PD=1.41536e-06 PS=1.44536e-06 $X=1500 $Y=660 $dt=0
M2 gnd3i! B Q gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.30162e-13 AS=2.28113e-13 PD=1.43036e-06 PS=1.41536e-06 $X=2340 $Y=660 $dt=0
M3 Q B gnd3i! gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=2.28113e-13 AS=2.30162e-13 PD=1.41536e-06 PS=1.43036e-06 $X=3230 $Y=660 $dt=0
M4 gnd3i! 7 Q gnd3i! ne3i L=3.4889e-07 W=9.00355e-07 AD=4.20212e-13 AS=2.28113e-13 PD=2.75536e-06 PS=1.41536e-06 $X=4070 $Y=660 $dt=0
M5 vdd3i! AN 7 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.998e-13 AS=6.768e-13 PD=2.595e-06 PS=3.78e-06 $X=620 $Y=2410 $dt=1
M6 9 7 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.115e-13 AS=6.998e-13 PD=1.71e-06 PS=2.595e-06 $X=1755 $Y=2410 $dt=1
M7 Q B 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.8775e-13 AS=2.115e-13 PD=1.96e-06 PS=1.71e-06 $X=2355 $Y=2410 $dt=1
M8 8 B Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.115e-13 AS=3.8775e-13 PD=1.71e-06 PS=1.96e-06 $X=3205 $Y=2410 $dt=1
M9 vdd3i! 7 8 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.3642e-12 AS=2.115e-13 PD=5.11e-06 PS=1.71e-06 $X=3805 $Y=2410 $dt=1
.ends NO2I1JI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX12                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX12 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=28
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=4.148e-13 AS=3.84e-13 PD=1.98e-06 PS=2.56e-06 $X=620 $Y=750 $dt=0
M1 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=4.148e-13 PD=1.34e-06 PS=1.98e-06 $X=1710 $Y=750 $dt=0
M2 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=2600 $Y=750 $dt=0
M3 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=3570 $Y=750 $dt=0
M4 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=4460 $Y=750 $dt=0
M5 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=5430 $Y=750 $dt=0
M6 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=6320 $Y=750 $dt=0
M7 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=7290 $Y=750 $dt=0
M8 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.404e-13 AS=2.16e-13 PD=1.86e-06 PS=1.34e-06 $X=8180 $Y=750 $dt=0
M9 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.16e-13 AS=3.404e-13 PD=1.34e-06 PS=1.86e-06 $X=9150 $Y=750 $dt=0
M10 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8e-07 AD=2.194e-13 AS=2.16e-13 PD=1.36e-06 PS=1.34e-06 $X=10040 $Y=750 $dt=0
M11 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.84e-13 AS=2.194e-13 PD=2.56e-06 PS=1.36e-06 $X=10930 $Y=750 $dt=0
M12 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=5.79287e-13 PD=1.86506e-06 PS=3.69506e-06 $X=475 $Y=2410 $dt=1
M13 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1315 $Y=2410 $dt=1
M14 6 A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=1865 $Y=2410 $dt=1
M15 vdd3i! A 6 vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=2705 $Y=2410 $dt=1
M16 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=3255 $Y=2410 $dt=1
M17 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=4095 $Y=2410 $dt=1
M18 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=4645 $Y=2410 $dt=1
M19 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=5485 $Y=2410 $dt=1
M20 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=6035 $Y=2410 $dt=1
M21 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=6875 $Y=2410 $dt=1
M22 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=7425 $Y=2410 $dt=1
M23 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=8265 $Y=2410 $dt=1
M24 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=8815 $Y=2410 $dt=1
M25 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.83187e-13 AS=2.54913e-13 PD=1.86506e-06 PS=1.86506e-06 $X=9655 $Y=2410 $dt=1
M26 Q 6 vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=2.83187e-13 PD=1.86506e-06 PS=1.86506e-06 $X=10205 $Y=2410 $dt=1
M27 vdd3i! 6 Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=8.53088e-13 AS=2.54913e-13 PD=4.55506e-06 PS=1.86506e-06 $X=11045 $Y=2410 $dt=1
.ends BUJI3VX12

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INJI3VX3                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INJI3VX3 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=5 EP=4 FDC=5
M0 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=7.586e-13 PD=1.43e-06 PS=3.76e-06 $X=780 $Y=660 $dt=0
M1 gnd3i! A Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=7.586e-13 AS=2.403e-13 PD=3.76e-06 PS=1.43e-06 $X=1670 $Y=660 $dt=0
M2 Q A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.54913e-13 AS=6.12287e-13 PD=1.86506e-06 PS=3.78506e-06 $X=490 $Y=2410 $dt=1
M3 vdd3i! A Q vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=2.86587e-13 AS=2.54913e-13 PD=1.88506e-06 PS=1.86506e-06 $X=1330 $Y=2410 $dt=1
M4 Q A vdd3i! vdd3i! pe3i L=3.00566e-07 W=1.47006e-06 AD=5.51013e-13 AS=2.86587e-13 PD=3.69506e-06 PS=1.88506e-06 $X=1880 $Y=2410 $dt=1
.ends INJI3VX3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA4JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA4JI3VX0 vdd3i! gnd3i! D Q C B A
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 11 D gnd3i! gnd3i! ne3i L=3.5e-07 W=8e-07 AD=1.2e-13 AS=7.868e-13 PD=1.1e-06 PS=3.82e-06 $X=810 $Y=750 $dt=0
M1 10 C 11 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=1.2e-13 AS=1.2e-13 PD=1.1e-06 PS=1.1e-06 $X=1460 $Y=750 $dt=0
M2 9 B 10 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=1.2e-13 AS=1.2e-13 PD=1.1e-06 PS=1.1e-06 $X=2110 $Y=750 $dt=0
M3 Q A 9 gnd3i! ne3i L=3.5e-07 W=8e-07 AD=3.84e-13 AS=1.2e-13 PD=2.56e-06 PS=1.1e-06 $X=2760 $Y=750 $dt=0
M4 Q D vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=9.882e-13 PD=1.24e-06 PS=3.92e-06 $X=540 $Y=2410 $dt=1
M5 vdd3i! C Q vdd3i! pe3i L=3e-07 W=7e-07 AD=9.882e-13 AS=1.89e-13 PD=3.92e-06 PS=1.24e-06 $X=1380 $Y=2410 $dt=1
M6 Q B vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=9.882e-13 PD=1.24e-06 PS=3.92e-06 $X=2240 $Y=2410 $dt=1
M7 vdd3i! A Q vdd3i! pe3i L=3e-07 W=7e-07 AD=9.882e-13 AS=1.89e-13 PD=3.92e-06 PS=1.24e-06 $X=3080 $Y=2410 $dt=1
.ends NA4JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OR3JI3VX1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OR3JI3VX1 vdd3i! gnd3i! A B C Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 gnd3i! A 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.482e-13 AS=2.016e-13 PD=2.04e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 8 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.116e-13 AS=2.482e-13 PD=1.78e-06 PS=2.04e-06 $X=1390 $Y=1310 $dt=0
M2 gnd3i! C 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.66689e-13 AS=2.116e-13 PD=1.17398e-06 PS=1.78e-06 $X=2160 $Y=1130 $dt=0
M3 Q 8 gnd3i! gnd3i! ne3i L=3.50112e-07 W=8.98284e-07 AD=4.174e-13 AS=3.56511e-13 PD=2.72828e-06 PS=2.51087e-06 $X=2970 $Y=660 $dt=0
M4 10 A 8 vdd3i! pe3i L=3e-07 W=1e-06 AD=1.375e-13 AS=4.8e-13 PD=1.275e-06 PS=2.96e-06 $X=670 $Y=2720 $dt=1
M5 9 B 10 vdd3i! pe3i L=3e-07 W=1e-06 AD=1.375e-13 AS=1.375e-13 PD=1.275e-06 PS=1.275e-06 $X=1245 $Y=2720 $dt=1
M6 vdd3i! C 9 vdd3i! pe3i L=3e-07 W=1e-06 AD=5.59502e-13 AS=1.375e-13 PD=2.19087e-06 PS=1.275e-06 $X=1820 $Y=2720 $dt=1
M7 Q 8 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=7.88898e-13 PD=3.78e-06 PS=3.08913e-06 $X=3000 $Y=2410 $dt=1
.ends OR3JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO3JI3VX1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO3JI3VX1 vdd3i! gnd3i! C Q B A
*.DEVICECLIMB
** N=9 EP=6 FDC=6
M0 Q C gnd3i! gnd3i! ne3i L=3.4986e-07 W=8.92071e-07 AD=2.37813e-13 AS=4.30337e-13 PD=1.42707e-06 PS=2.76707e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! B Q gnd3i! ne3i L=3.4986e-07 W=8.92071e-07 AD=2.40287e-13 AS=2.37813e-13 PD=1.44207e-06 PS=1.42707e-06 $X=1500 $Y=660 $dt=0
M2 Q A gnd3i! gnd3i! ne3i L=3.4986e-07 W=8.92071e-07 AD=4.29162e-13 AS=2.40287e-13 PD=2.74707e-06 PS=1.44207e-06 $X=2390 $Y=660 $dt=0
M3 9 C vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=1.3994e-12 PD=1.72e-06 PS=5.15e-06 $X=955 $Y=2410 $dt=1
M4 8 B 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=2.1855e-13 PD=1.72e-06 PS=1.72e-06 $X=1565 $Y=2410 $dt=1
M5 Q A 8 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=2.1855e-13 PD=3.78e-06 PS=1.72e-06 $X=2175 $Y=2410 $dt=1
.ends NO3JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: FAJI3VX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt FAJI3VX1 vdd3i! gnd3i! S CI B A CO
*.DEVICECLIMB
** N=20 EP=7 FDC=28
M0 gnd3i! 12 S gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.361e-13 AS=4.272e-13 PD=2.76e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 15 CI 12 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=7.375e-14 AS=2.832e-13 PD=8.4e-07 PS=2.14e-06 $X=2220 $Y=960 $dt=0
M2 14 B 15 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=7.375e-14 AS=7.375e-14 PD=8.4e-07 PS=8.4e-07 $X=2820 $Y=960 $dt=0
M3 gnd3i! A 14 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=2.34033e-13 AS=7.375e-14 PD=1.52158e-06 PS=8.4e-07 $X=3420 $Y=960 $dt=0
M4 13 CI gnd3i! gnd3i! ne3i L=3.5e-07 W=5.5e-07 AD=1.485e-13 AS=2.18167e-13 PD=1.09e-06 PS=1.41842e-06 $X=4350 $Y=660 $dt=0
M5 gnd3i! A 13 gnd3i! ne3i L=3.5e-07 W=5.5e-07 AD=2.5017e-13 AS=1.485e-13 PD=1.58058e-06 PS=1.09e-06 $X=5240 $Y=660 $dt=0
M6 13 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=1.296e-13 AS=2.1833e-13 PD=1.02e-06 PS=1.37942e-06 $X=6220 $Y=960 $dt=0
M7 12 10 13 gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=2.304e-13 AS=1.296e-13 PD=1.92e-06 PS=1.02e-06 $X=7110 $Y=960 $dt=0
M8 gnd3i! 10 CO gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=3.345e-13 AS=2.832e-13 PD=1.73e-06 PS=2.14e-06 $X=8700 $Y=960 $dt=0
M9 11 A gnd3i! gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=7.375e-14 AS=3.345e-13 PD=8.4e-07 PS=1.73e-06 $X=9830 $Y=960 $dt=0
M10 10 B 11 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=1.593e-13 AS=7.375e-14 PD=1.13e-06 PS=8.4e-07 $X=10430 $Y=960 $dt=0
M11 9 CI 10 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=1.593e-13 AS=1.593e-13 PD=1.13e-06 PS=1.13e-06 $X=11320 $Y=960 $dt=0
M12 gnd3i! B 9 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=4.382e-13 AS=1.593e-13 PD=1.95e-06 PS=1.13e-06 $X=12210 $Y=960 $dt=0
M13 9 A gnd3i! gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=3.068e-13 AS=4.382e-13 PD=2.22e-06 PS=1.95e-06 $X=13550 $Y=960 $dt=0
M14 vdd3i! 12 S vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.6395e-13 AS=7.1205e-13 PD=4.52213e-06 PS=3.83e-06 $X=645 $Y=2410 $dt=1
M15 vdd3i! CI 17 vdd3i! pe3i L=3e-07 W=1.03e-06 AD=4.8155e-13 AS=4.79437e-13 PD=2.35e-06 PS=3.03778e-06 $X=2125 $Y=2490 $dt=1
M16 17 B vdd3i! vdd3i! pe3i L=3e-07 W=1.03e-06 AD=3.0385e-13 AS=4.8155e-13 PD=1.62e-06 PS=2.35e-06 $X=3095 $Y=2490 $dt=1
M17 vdd3i! A 17 vdd3i! pe3i L=3e-07 W=1.03e-06 AD=4.1015e-13 AS=3.0385e-13 PD=2.01e-06 PS=1.62e-06 $X=3985 $Y=2490 $dt=1
M18 20 A vdd3i! vdd3i! pe3i L=3e-07 W=1.03e-06 AD=1.545e-13 AS=4.1015e-13 PD=1.33e-06 PS=2.01e-06 $X=4955 $Y=2490 $dt=1
M19 19 B 20 vdd3i! pe3i L=3e-07 W=1.03e-06 AD=1.545e-13 AS=1.545e-13 PD=1.33e-06 PS=1.33e-06 $X=5555 $Y=2490 $dt=1
M20 12 CI 19 vdd3i! pe3i L=3e-07 W=1.03e-06 AD=3.0385e-13 AS=1.545e-13 PD=1.62e-06 PS=1.33e-06 $X=6155 $Y=2490 $dt=1
M21 17 10 12 vdd3i! pe3i L=3e-07 W=1.03e-06 AD=6.9155e-13 AS=3.0385e-13 PD=3.77e-06 PS=1.62e-06 $X=7045 $Y=2490 $dt=1
M22 vdd3i! 10 CO vdd3i! pe3i L=3e-07 W=1.11e-06 AD=4.54624e-13 AS=5.6055e-13 PD=2.27286e-06 PS=3.23e-06 $X=8675 $Y=2410 $dt=1
M23 16 A vdd3i! vdd3i! pe3i L=3e-07 W=9.9e-07 AD=2.9205e-13 AS=4.05476e-13 PD=1.58e-06 PS=2.02714e-06 $X=9645 $Y=2530 $dt=1
M24 vdd3i! B 16 vdd3i! pe3i L=3e-07 W=9.9e-07 AD=5.763e-13 AS=2.9205e-13 PD=3.59e-06 PS=1.58e-06 $X=10535 $Y=2530 $dt=1
M25 10 CI 16 vdd3i! pe3i L=3e-07 W=1e-06 AD=2.95e-13 AS=4.65e-13 PD=1.59e-06 PS=3.01e-06 $X=12085 $Y=2520 $dt=1
M26 18 B 10 vdd3i! pe3i L=3e-07 W=1e-06 AD=1.5e-13 AS=2.95e-13 PD=1.3e-06 PS=1.59e-06 $X=12975 $Y=2520 $dt=1
M27 vdd3i! A 18 vdd3i! pe3i L=3e-07 W=1e-06 AD=8.18e-13 AS=1.5e-13 PD=4.39e-06 PS=1.3e-06 $X=13575 $Y=2520 $dt=1
.ends FAJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX4                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX4 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=11
M0 6 A gnd3i! gnd3i! ne3i L=3.5e-07 W=5.95e-07 AD=1.6065e-13 AS=5.803e-13 PD=1.135e-06 PS=3.52e-06 $X=660 $Y=955 $dt=0
M1 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=5.95e-07 AD=3.92379e-13 AS=1.6065e-13 PD=1.69084e-06 PS=1.135e-06 $X=1550 $Y=955 $dt=0
M2 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=5.86921e-13 PD=1.43e-06 PS=2.52916e-06 $X=2770 $Y=660 $dt=0
M3 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=3660 $Y=660 $dt=0
M4 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=3.494e-13 PD=2.74e-06 PS=1.86e-06 $X=4630 $Y=660 $dt=0
M5 6 A vdd3i! vdd3i! pe3i L=3e-07 W=1.1e-06 AD=2.97e-13 AS=9.042e-13 PD=1.64e-06 PS=4.66e-06 $X=710 $Y=2410 $dt=1
M6 vdd3i! A 6 vdd3i! pe3i L=3e-07 W=1.1e-06 AD=4.45401e-13 AS=2.97e-13 PD=2.09699e-06 PS=1.64e-06 $X=1550 $Y=2410 $dt=1
M7 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=5.91049e-13 PD=1.87971e-06 PS=2.78272e-06 $X=2445 $Y=2410 $dt=1
M8 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=3.3675e-13 AS=2.751e-13 PD=1.92971e-06 PS=1.87971e-06 $X=3285 $Y=2410 $dt=1
M9 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=3.3675e-13 PD=1.87971e-06 PS=1.92971e-06 $X=3935 $Y=2410 $dt=1
M10 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=6.3285e-13 AS=2.751e-13 PD=3.75971e-06 PS=1.87971e-06 $X=4775 $Y=2410 $dt=1
.ends BUJI3VX4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INJI3VX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INJI3VX1 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=5 EP=4 FDC=2
M0 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=6e-07 AD=2.88e-13 AS=6.428e-13 PD=2.16e-06 PS=3.62e-06 $X=710 $Y=950 $dt=0
M1 Q A vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=1.0562e-12 PD=3.78e-06 PS=4.76e-06 $X=760 $Y=2410 $dt=1
.ends INJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DLY2JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DLY2JI3VX1 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=12 EP=4 FDC=12
M0 gnd3i! A 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=3.577e-13 AS=2.016e-13 PD=1.79e-06 PS=1.8e-06 $X=620 $Y=660 $dt=0
M1 8 10 gnd3i! gnd3i! ne3i L=8e-07 W=4.2e-07 AD=2.548e-13 AS=3.577e-13 PD=1.7e-06 PS=1.79e-06 $X=1990 $Y=660 $dt=0
M2 8 10 9 gnd3i! ne3i L=8e-07 W=4.2e-07 AD=2.548e-13 AS=2.016e-13 PD=1.7e-06 PS=1.8e-06 $X=1990 $Y=1360 $dt=0
M3 gnd3i! 9 7 gnd3i! ne3i L=1e-06 W=4.2e-07 AD=3.42444e-13 AS=2.1e-13 PD=1.66718e-06 PS=1.62e-06 $X=3950 $Y=660 $dt=0
M4 6 9 7 gnd3i! ne3i L=1e-06 W=4.2e-07 AD=2.10588e-13 AS=2.1e-13 PD=1.81778e-06 PS=1.62e-06 $X=3950 $Y=1360 $dt=0
M5 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=7.25656e-13 PD=2.74e-06 PS=3.53282e-06 $X=6310 $Y=660 $dt=0
M6 vdd3i! A 10 vdd3i! pe3i L=3e-07 W=7e-07 AD=5.42937e-13 AS=3.535e-13 PD=2.69375e-06 PS=2.41e-06 $X=645 $Y=3120 $dt=1
M7 12 10 9 vdd3i! pe3i L=7.4e-07 W=4.2e-07 AD=2.8095e-13 AS=2.0035e-13 PD=1.785e-06 PS=1.77071e-06 $X=2050 $Y=2640 $dt=1
M8 12 10 vdd3i! vdd3i! pe3i L=7.4e-07 W=4.2e-07 AD=2.8095e-13 AS=3.25762e-13 PD=1.785e-06 PS=1.61625e-06 $X=2050 $Y=3400 $dt=1
M9 6 9 11 vdd3i! pe3i L=1e-06 W=4.2e-07 AD=2.856e-13 AS=2.479e-13 PD=2.2e-06 PS=1.715e-06 $X=4030 $Y=2660 $dt=1
M10 vdd3i! 9 11 vdd3i! pe3i L=1e-06 W=4.2e-07 AD=2.62018e-13 AS=2.479e-13 PD=1.40689e-06 PS=1.715e-06 $X=4030 $Y=3400 $dt=1
M11 Q 6 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=7.1205e-13 AS=8.79632e-13 PD=3.83e-06 PS=4.72311e-06 $X=6335 $Y=2410 $dt=1
.ends DLY2JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: SDFRRQJI3VX1                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt SDFRRQJI3VX1 vdd3i! gnd3i! SE SD RN D C Q
*.DEVICECLIMB
** N=31 EP=8 FDC=39
M0 gnd3i! SE 25 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.11575e-13 AS=2.016e-13 PD=1.6275e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 13 RN gnd3i! gnd3i! ne3i L=3.5e-07 W=5.4e-07 AD=2.079e-13 AS=2.72025e-13 PD=1.4625e-06 PS=2.0925e-06 $X=1410 $Y=660 $dt=0
M2 24 SE 13 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.617e-13 PD=6.7e-07 PS=1.1375e-06 $X=2340 $Y=960 $dt=0
M3 12 SD 24 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.163e-13 AS=5.25e-14 PD=1.45e-06 PS=6.7e-07 $X=2940 $Y=960 $dt=0
M4 23 D 12 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.163e-13 PD=6.7e-07 PS=1.45e-06 $X=3910 $Y=1000 $dt=0
M5 13 25 23 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=5.25e-14 PD=1.8e-06 PS=6.7e-07 $X=4510 $Y=1000 $dt=0
M6 gnd3i! 20 22 gnd3i! ne3i L=3.5e-07 W=7.2e-07 AD=3.01862e-13 AS=3.456e-13 PD=1.65084e-06 PS=2.4e-06 $X=6100 $Y=1090 $dt=0
M7 11 RN gnd3i! gnd3i! ne3i L=3.5e-07 W=8.85e-07 AD=2.20538e-13 AS=3.71038e-13 PD=1.77e-06 PS=2.02916e-06 $X=7070 $Y=925 $dt=0
M8 21 22 11 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.04662e-13 PD=6.7e-07 PS=8.4e-07 $X=7840 $Y=1390 $dt=0
M9 20 18 21 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=8440 $Y=1390 $dt=0
M10 12 19 20 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=1.134e-13 PD=1.8e-06 PS=9.6e-07 $X=9330 $Y=1390 $dt=0
M11 gnd3i! C 19 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.722e-13 AS=2.016e-13 PD=1.24e-06 PS=1.8e-06 $X=10920 $Y=1390 $dt=0
M12 18 19 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=1.722e-13 PD=1.8e-06 PS=1.24e-06 $X=11930 $Y=1390 $dt=0
M13 17 22 10 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.016e-13 PD=6.7e-07 PS=1.8e-06 $X=13520 $Y=1020 $dt=0
M14 16 18 17 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.25e-14 PD=9.6e-07 PS=6.7e-07 $X=14120 $Y=1020 $dt=0
M15 15 19 16 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=1.134e-13 PD=6.7e-07 PS=9.6e-07 $X=15010 $Y=1020 $dt=0
M16 10 14 15 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.47785e-13 AS=5.25e-14 PD=9.42595e-07 PS=6.7e-07 $X=15610 $Y=1020 $dt=0
M17 gnd3i! RN 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.9815e-13 AS=3.13165e-13 PD=1.56e-06 PS=1.9974e-06 $X=16540 $Y=660 $dt=0
M18 14 16 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=2.9815e-13 PD=2.74e-06 PS=1.56e-06 $X=17560 $Y=660 $dt=0
M19 Q 16 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=6.098e-13 PD=2.74e-06 PS=3.52e-06 $X=19190 $Y=660 $dt=0
M20 vdd3i! SE 25 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=5.776e-13 AS=3.456e-13 PD=2.10667e-06 PS=2.4e-06 $X=620 $Y=2800 $dt=1
M21 31 25 vdd3i! vdd3i! pe3i L=3e-07 W=9e-07 AD=1.125e-13 AS=7.22e-13 PD=1.15e-06 PS=2.63333e-06 $X=2030 $Y=2620 $dt=1
M22 28 SD 31 vdd3i! pe3i L=3e-07 W=9e-07 AD=2.43e-13 AS=1.125e-13 PD=1.44e-06 PS=1.15e-06 $X=2580 $Y=2620 $dt=1
M23 30 D 28 vdd3i! pe3i L=3e-07 W=9e-07 AD=1.125e-13 AS=2.43e-13 PD=1.15e-06 PS=1.44e-06 $X=3420 $Y=2620 $dt=1
M24 vdd3i! SE 30 vdd3i! pe3i L=3e-07 W=9e-07 AD=3.80558e-13 AS=1.125e-13 PD=1.98274e-06 PS=1.15e-06 $X=3970 $Y=2620 $dt=1
M25 22 20 vdd3i! vdd3i! pe3i L=3e-07 W=1.07e-06 AD=5.136e-13 AS=4.52442e-13 PD=3.1e-06 PS=2.35726e-06 $X=4890 $Y=2745 $dt=1
M26 vdd3i! RN 20 vdd3i! pe3i L=3e-07 W=1.02e-06 AD=9.30148e-13 AS=4.896e-13 PD=3.58417e-06 PS=3e-06 $X=6430 $Y=2800 $dt=1
M27 29 22 vdd3i! vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=3.83002e-13 PD=6.7e-07 PS=1.47583e-06 $X=7890 $Y=3060 $dt=1
M28 20 19 29 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=1.218e-13 AS=5.25e-14 PD=9.22677e-07 PS=6.7e-07 $X=8440 $Y=3060 $dt=1
M29 28 18 20 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.08e-13 AS=2.465e-13 PD=2.66e-06 PS=1.86732e-06 $X=9285 $Y=2670 $dt=1
M30 19 C vdd3i! vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.0675e-13 AS=6.327e-13 PD=2.37071e-06 PS=3.56e-06 $X=10970 $Y=2735 $dt=1
M31 vdd3i! 19 18 vdd3i! pe3i L=3e-07 W=7.2e-07 AD=3.27981e-13 AS=4.01587e-13 PD=1.59258e-06 PS=3.03778e-06 $X=12390 $Y=2800 $dt=1
M32 27 22 vdd3i! vdd3i! pe3i L=3e-07 W=7.9e-07 AD=1.16525e-13 AS=3.59869e-13 PD=1.085e-06 PS=1.74742e-06 $X=13570 $Y=2730 $dt=1
M33 16 19 27 vdd3i! pe3i L=3e-07 W=7.9e-07 AD=2.25379e-13 AS=1.16525e-13 PD=1.73669e-06 PS=1.085e-06 $X=14165 $Y=2730 $dt=1
M34 26 18 16 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=5.25e-14 AS=1.19821e-13 PD=6.7e-07 PS=9.23306e-07 $X=15005 $Y=3100 $dt=1
M35 vdd3i! 14 26 vdd3i! pe3i L=3e-07 W=4.2e-07 AD=6.29844e-13 AS=5.25e-14 PD=2.86017e-06 PS=6.7e-07 $X=15555 $Y=3100 $dt=1
M36 vdd3i! RN 16 vdd3i! pe3i L=3e-07 W=7.9e-07 AD=1.18471e-12 AS=3.19387e-13 PD=5.37983e-06 PS=2.5195e-06 $X=16775 $Y=2410 $dt=1
M37 vdd3i! 16 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=6.768e-13 PD=1.95e-06 PS=3.78e-06 $X=18400 $Y=2410 $dt=1
M38 Q 16 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=3.807e-13 PD=3.78e-06 PS=1.95e-06 $X=19240 $Y=2410 $dt=1
.ends SDFRRQJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: BUJI3VX3                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt BUJI3VX3 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=6 EP=4 FDC=7
M0 gnd3i! A 6 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=5.23e-13 AS=4.272e-13 PD=2.14e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 Q 6 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.5365e-13 AS=5.23e-13 PD=1.46e-06 PS=2.14e-06 $X=1870 $Y=660 $dt=0
M2 gnd3i! 6 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=7.586e-13 AS=2.5365e-13 PD=3.76e-06 PS=1.46e-06 $X=2790 $Y=660 $dt=0
M3 vdd3i! A 6 vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=6.11825e-13 AS=5.712e-13 PD=2.51971e-06 PS=3.70971e-06 $X=620 $Y=2410 $dt=1
M4 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=6.11825e-13 PD=1.87971e-06 PS=2.51971e-06 $X=1510 $Y=2410 $dt=1
M5 vdd3i! 6 Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=3.3675e-13 AS=2.751e-13 PD=1.92971e-06 PS=1.87971e-06 $X=2350 $Y=2410 $dt=1
M6 Q 6 vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=5.712e-13 AS=3.3675e-13 PD=3.70971e-06 PS=1.92971e-06 $X=3000 $Y=2410 $dt=1
.ends BUJI3VX3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INJI3VX0                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INJI3VX0 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=5 EP=4 FDC=2
M0 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=6.248e-13 PD=1.8e-06 PS=3.62e-06 $X=710 $Y=1130 $dt=0
M1 Q A vdd3i! vdd3i! pe3i L=3e-07 W=9.4e-07 AD=4.512e-13 AS=1.0092e-12 PD=2.84e-06 PS=4.76e-06 $X=760 $Y=2410 $dt=1
.ends INJI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA2JI3VX0 vdd3i! gnd3i! B Q A
*.DEVICECLIMB
** N=7 EP=5 FDC=4
M0 7 B gnd3i! gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=5.892e-13 PD=8.1e-07 PS=3.54e-06 $X=670 $Y=990 $dt=0
M1 Q A 7 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=2.688e-13 AS=7e-14 PD=2.08e-06 PS=8.1e-07 $X=1270 $Y=990 $dt=0
M2 Q B vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=1.1114e-12 PD=1.24e-06 PS=4.94e-06 $X=550 $Y=2410 $dt=1
M3 vdd3i! A Q vdd3i! pe3i L=3e-07 W=7e-07 AD=1.1114e-12 AS=1.89e-13 PD=4.94e-06 PS=1.24e-06 $X=1390 $Y=2410 $dt=1
.ends NA2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AO22JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AO22JI3VX1 vdd3i! gnd3i! B A C D Q
*.DEVICECLIMB
** N=12 EP=7 FDC=10
M0 11 B gnd3i! gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=5.768e-13 PD=8.1e-07 PS=3.52e-06 $X=660 $Y=990 $dt=0
M1 10 A 11 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=1.68e-13 AS=7e-14 PD=1.16e-06 PS=8.1e-07 $X=1260 $Y=990 $dt=0
M2 9 C 10 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=1.68e-13 PD=8.1e-07 PS=1.16e-06 $X=2210 $Y=990 $dt=0
M3 gnd3i! D 9 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=3.96017e-13 AS=7e-14 PD=1.66069e-06 PS=8.1e-07 $X=2810 $Y=990 $dt=0
M4 Q 10 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=6.29383e-13 PD=2.74e-06 PS=2.63931e-06 $X=4070 $Y=660 $dt=0
M5 vdd3i! B 12 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=2.295e-13 AS=4.868e-13 PD=1.39e-06 PS=3.75e-06 $X=460 $Y=2490 $dt=1
M6 12 A vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.868e-13 AS=2.295e-13 PD=3.75e-06 PS=1.39e-06 $X=1300 $Y=2490 $dt=1
M7 10 C 12 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=2.295e-13 AS=4.868e-13 PD=1.39e-06 PS=3.75e-06 $X=2020 $Y=2490 $dt=1
M8 12 D 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.868e-13 AS=2.295e-13 PD=3.75e-06 PS=1.39e-06 $X=2860 $Y=2490 $dt=1
M9 Q 10 vdd3i! vdd3i! pe3i L=3.01705e-07 W=1.47627e-06 AD=5.312e-13 AS=7.778e-13 PD=3.68627e-06 PS=4.46627e-06 $X=4120 $Y=2410 $dt=1
.ends AO22JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OR4JI3VX2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OR4JI3VX2 vdd3i! gnd3i! C D Q B A
*.DEVICECLIMB
** N=14 EP=7 FDC=16
M0 10 C gnd3i! gnd3i! ne3i L=3.5e-07 W=7e-07 AD=1.9155e-13 AS=3.417e-13 PD=1.255e-06 PS=2.39e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! D 10 gnd3i! ne3i L=3.5e-07 W=7e-07 AD=2.07711e-13 AS=1.9155e-13 PD=1.27673e-06 PS=1.255e-06 $X=1510 $Y=660 $dt=0
M2 12 10 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=2.64089e-13 PD=1.14e-06 PS=1.62327e-06 $X=2420 $Y=660 $dt=0
M3 Q 9 12 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=1.1125e-13 PD=1.43e-06 PS=1.14e-06 $X=3020 $Y=660 $dt=0
M4 11 9 Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.2015e-13 AS=2.403e-13 PD=1.16e-06 PS=1.43e-06 $X=3910 $Y=660 $dt=0
M5 gnd3i! 10 11 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.54126e-13 AS=1.2015e-13 PD=1.60088e-06 PS=1.16e-06 $X=4530 $Y=660 $dt=0
M6 9 B gnd3i! gnd3i! ne3i L=3.5e-07 W=7e-07 AD=1.9155e-13 AS=1.99874e-13 PD=1.255e-06 PS=1.25912e-06 $X=5420 $Y=660 $dt=0
M7 gnd3i! A 9 gnd3i! ne3i L=3.5e-07 W=7e-07 AD=3.417e-13 AS=1.9155e-13 PD=2.39e-06 PS=1.255e-06 $X=6310 $Y=660 $dt=0
M8 14 C 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=6.768e-13 PD=1.66e-06 PS=3.78e-06 $X=710 $Y=2410 $dt=1
M9 vdd3i! D 14 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=5.47043e-13 AS=1.7625e-13 PD=2.41704e-06 PS=1.66e-06 $X=1260 $Y=2410 $dt=1
M10 Q 10 vdd3i! vdd3i! pe3i L=2.99799e-07 W=1.41828e-06 AD=3.622e-13 AS=5.50257e-13 PD=1.93828e-06 PS=2.43124e-06 $X=2210 $Y=2410 $dt=1
M11 vdd3i! 9 Q vdd3i! pe3i L=2.99799e-07 W=1.41828e-06 AD=4.987e-13 AS=3.622e-13 PD=2.36828e-06 PS=1.93828e-06 $X=3050 $Y=2410 $dt=1
M12 Q 9 vdd3i! vdd3i! pe3i L=2.99799e-07 W=1.41828e-06 AD=3.622e-13 AS=4.987e-13 PD=1.93828e-06 PS=2.36828e-06 $X=3930 $Y=2410 $dt=1
M13 vdd3i! 10 Q vdd3i! pe3i L=2.99799e-07 W=1.41828e-06 AD=5.8556e-13 AS=3.622e-13 PD=2.47136e-06 PS=1.93828e-06 $X=4770 $Y=2410 $dt=1
M14 13 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=5.8214e-13 PD=1.66e-06 PS=2.45692e-06 $X=5760 $Y=2410 $dt=1
M15 9 A 13 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=1.7625e-13 PD=3.78e-06 PS=1.66e-06 $X=6310 $Y=2410 $dt=1
.ends OR4JI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INJI3VX2                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INJI3VX2 vdd3i! gnd3i! A Q
*.DEVICECLIMB
** N=5 EP=4 FDC=4
M0 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=1.296e-13 AS=4.408e-13 PD=1.02e-06 PS=3.52e-06 $X=500 $Y=1070 $dt=0
M1 gnd3i! A Q gnd3i! ne3i L=3.5e-07 W=4.8e-07 AD=4.408e-13 AS=1.296e-13 PD=3.52e-06 PS=1.02e-06 $X=1390 $Y=1070 $dt=0
M2 Q A vdd3i! vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=2.751e-13 AS=8.151e-13 PD=1.87971e-06 PS=4.50971e-06 $X=560 $Y=2410 $dt=1
M3 vdd3i! A Q vdd3i! pe3i L=3.00472e-07 W=1.45971e-06 AD=8.01e-13 AS=2.751e-13 PD=4.48971e-06 PS=1.87971e-06 $X=1400 $Y=2410 $dt=1
.ends INJI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AO21JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AO21JI3VX1 vdd3i! gnd3i! B A C Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 9 B gnd3i! gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=5.768e-13 PD=8.1e-07 PS=3.52e-06 $X=660 $Y=990 $dt=0
M1 8 A 9 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=1.708e-13 AS=7e-14 PD=1.17e-06 PS=8.1e-07 $X=1260 $Y=990 $dt=0
M2 gnd3i! C 8 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=3.94626e-13 AS=1.708e-13 PD=1.68386e-06 PS=1.17e-06 $X=2220 $Y=990 $dt=0
M3 Q 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=6.27174e-13 PD=2.74e-06 PS=2.67614e-06 $X=3510 $Y=660 $dt=0
M4 vdd3i! B 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=3.8185e-13 AS=4.08e-13 PD=2.53e-06 PS=2.66e-06 $X=620 $Y=2410 $dt=1
M5 10 A vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=2.295e-13 AS=3.8185e-13 PD=1.39e-06 PS=2.53e-06 $X=1340 $Y=2410 $dt=1
M6 8 C 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.08e-13 AS=2.295e-13 PD=2.66e-06 PS=1.39e-06 $X=2180 $Y=2410 $dt=1
M7 Q 8 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=7.0775e-13 PD=3.78e-06 PS=4.73e-06 $X=3560 $Y=2410 $dt=1
.ends AO21JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO2I1JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO2I1JI3VX1 vdd3i! gnd3i! AN Q B
*.DEVICECLIMB
** N=8 EP=5 FDC=6
M0 gnd3i! AN 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.78131e-13 AS=2.016e-13 PD=1.19267e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 Q 7 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.4285e-13 AS=3.77469e-13 PD=1.445e-06 PS=2.52733e-06 $X=1460 $Y=660 $dt=0
M2 gnd3i! B Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=6.098e-13 AS=2.4285e-13 PD=3.52e-06 PS=1.445e-06 $X=2350 $Y=660 $dt=0
M3 vdd3i! AN 7 vdd3i! pe3i L=3e-07 W=7e-07 AD=4.32009e-13 AS=3.36e-13 PD=1.71185e-06 PS=2.36e-06 $X=620 $Y=2410 $dt=1
M4 8 7 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=8.70191e-13 PD=1.66e-06 PS=3.44815e-06 $X=1740 $Y=2410 $dt=1
M5 Q B 8 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=1.7625e-13 PD=3.78e-06 PS=1.66e-06 $X=2290 $Y=2410 $dt=1
.ends NO2I1JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA3JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA3JI3VX0 vdd3i! gnd3i! C Q B A
*.DEVICECLIMB
** N=9 EP=6 FDC=6
M0 9 C gnd3i! gnd3i! ne3i L=3.5e-07 W=7e-07 AD=8.75e-14 AS=5.605e-13 PD=9.5e-07 PS=3.52e-06 $X=630 $Y=850 $dt=0
M1 8 B 9 gnd3i! ne3i L=3.5e-07 W=7e-07 AD=8.75e-14 AS=8.75e-14 PD=9.5e-07 PS=9.5e-07 $X=1230 $Y=850 $dt=0
M2 Q A 8 gnd3i! ne3i L=3.5e-07 W=7e-07 AD=3.36e-13 AS=8.75e-14 PD=2.36e-06 PS=9.5e-07 $X=1830 $Y=850 $dt=0
M3 Q C vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=5.76467e-13 PD=1.24e-06 PS=3.21333e-06 $X=470 $Y=2580 $dt=1
M4 vdd3i! B Q vdd3i! pe3i L=3e-07 W=7e-07 AD=5.76467e-13 AS=1.89e-13 PD=3.21333e-06 PS=1.24e-06 $X=1310 $Y=2580 $dt=1
M5 Q A vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=4.708e-13 AS=5.76467e-13 PD=3.92e-06 PS=3.21333e-06 $X=2040 $Y=2470 $dt=1
.ends NA3JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OR2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OR2JI3VX0 vdd3i! gnd3i! A B Q
*.DEVICECLIMB
** N=8 EP=5 FDC=6
M0 7 A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.75467e-13 PD=9.6e-07 PS=2.95333e-06 $X=530 $Y=1130 $dt=0
M1 gnd3i! B 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.75467e-13 AS=1.134e-13 PD=2.95333e-06 PS=9.6e-07 $X=1420 $Y=1130 $dt=0
M2 Q 7 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=5.75467e-13 PD=1.8e-06 PS=2.95333e-06 $X=2390 $Y=1130 $dt=0
M3 8 A 7 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=4.08e-13 PD=1.1e-06 PS=2.66e-06 $X=620 $Y=2410 $dt=1
M4 vdd3i! B 8 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=8.28174e-13 AS=1.0625e-13 PD=2.99419e-06 PS=1.1e-06 $X=1170 $Y=2410 $dt=1
M5 Q 7 vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=3.36e-13 AS=6.82026e-13 PD=2.36e-06 PS=2.46581e-06 $X=2440 $Y=2410 $dt=1
.ends OR2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AO211JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AO211JI3VX1 vdd3i! gnd3i! B A C D Q
*.DEVICECLIMB
** N=12 EP=7 FDC=10
M0 10 B gnd3i! gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=5.768e-13 PD=8.1e-07 PS=3.52e-06 $X=660 $Y=990 $dt=0
M1 9 A 10 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=1.68e-13 AS=7e-14 PD=1.16e-06 PS=8.1e-07 $X=1260 $Y=990 $dt=0
M2 gnd3i! C 9 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=3.164e-13 AS=1.68e-13 PD=1.86e-06 PS=1.16e-06 $X=2210 $Y=990 $dt=0
M3 9 D gnd3i! gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=2.464e-13 AS=3.164e-13 PD=2.08e-06 PS=1.86e-06 $X=3180 $Y=990 $dt=0
M4 Q 9 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=5.0945e-13 PD=2.74e-06 PS=3.7e-06 $X=4630 $Y=660 $dt=0
M5 vdd3i! B 12 vdd3i! pe3i L=3e-07 W=1e-06 AD=4.168e-13 AS=4.8e-13 PD=2.53e-06 PS=2.96e-06 $X=620 $Y=2410 $dt=1
M6 12 A vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.95e-13 AS=4.168e-13 PD=1.59e-06 PS=2.53e-06 $X=1410 $Y=2410 $dt=1
M7 11 C 12 vdd3i! pe3i L=3e-07 W=1e-06 AD=1.5e-13 AS=2.95e-13 PD=1.3e-06 PS=1.59e-06 $X=2300 $Y=2410 $dt=1
M8 9 D 11 vdd3i! pe3i L=3e-07 W=1e-06 AD=4.66e-13 AS=1.5e-13 PD=3.28e-06 PS=1.3e-06 $X=2900 $Y=2410 $dt=1
M9 Q 9 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=1.01495e-12 PD=3.78e-06 PS=4.82e-06 $X=4680 $Y=2410 $dt=1
.ends AO211JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: HAJI3VX1                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt HAJI3VX1 vdd3i! gnd3i! S B A CO
*.DEVICECLIMB
** N=12 EP=6 FDC=14
M0 gnd3i! 8 S gnd3i! ne3i L=3.49889e-07 W=8.98284e-07 AD=4.998e-13 AS=4.174e-13 PD=3.41456e-06 PS=2.72828e-06 $X=600 $Y=660 $dt=0
M1 gnd3i! A 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.52e-13 PD=1.43e-06 PS=2.74e-06 $X=2070 $Y=660 $dt=0
M2 9 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.70969e-13 AS=2.403e-13 PD=1.71986e-06 PS=1.43e-06 $X=2960 $Y=660 $dt=0
M3 8 10 9 gnd3i! ne3i L=3.5e-07 W=5.9e-07 AD=3.632e-13 AS=1.79631e-13 PD=2.84284e-06 PS=1.14014e-06 $X=3850 $Y=960 $dt=0
M4 gnd3i! 10 CO gnd3i! ne3i L=3.5e-07 W=5.5e-07 AD=1.56292e-13 AS=2.4195e-13 PD=1.09236e-06 PS=2.03071e-06 $X=5380 $Y=1000 $dt=0
M5 11 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=2.52908e-13 PD=1.14e-06 PS=1.76764e-06 $X=6270 $Y=660 $dt=0
M6 10 A 11 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=1.1125e-13 PD=2.74e-06 PS=1.14e-06 $X=6870 $Y=660 $dt=0
M7 vdd3i! 8 S vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.07833e-13 AS=7.1205e-13 PD=2.97939e-06 PS=3.83e-06 $X=645 $Y=2410 $dt=1
M8 12 A vdd3i! vdd3i! pe3i L=3e-07 W=8.9e-07 AD=1.335e-13 AS=3.83667e-13 PD=1.19e-06 PS=1.88061e-06 $X=1615 $Y=2630 $dt=1
M9 8 B 12 vdd3i! pe3i L=3e-07 W=8.9e-07 AD=4.9565e-13 AS=1.335e-13 PD=2.12e-06 PS=1.19e-06 $X=2215 $Y=2630 $dt=1
M10 vdd3i! 10 8 vdd3i! pe3i L=3e-07 W=8.9e-07 AD=4.8925e-13 AS=4.9565e-13 PD=3.49e-06 PS=2.12e-06 $X=3525 $Y=2630 $dt=1
M11 vdd3i! 10 CO vdd3i! pe3i L=3e-07 W=1.11e-06 AD=4.3695e-13 AS=4.7415e-13 PD=2.09e-06 PS=3.23e-06 $X=4995 $Y=2410 $dt=1
M12 10 B vdd3i! vdd3i! pe3i L=3e-07 W=1.11e-06 AD=3.2745e-13 AS=4.3695e-13 PD=1.7e-06 PS=2.09e-06 $X=5965 $Y=2410 $dt=1
M13 vdd3i! A 10 vdd3i! pe3i L=3e-07 W=1.11e-06 AD=8.7795e-13 AS=3.2745e-13 PD=4.61e-06 PS=1.7e-06 $X=6855 $Y=2410 $dt=1
.ends HAJI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OA21JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OA21JI3VX1 vdd3i! gnd3i! C A B Q
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 8 C 9 gnd3i! ne3i L=3.5e-07 W=5.4e-07 AD=3.313e-13 AS=2.97e-13 PD=1.95333e-06 PS=2.18e-06 $X=690 $Y=660 $dt=0
M1 8 A gnd3i! gnd3i! ne3i L=3.5e-07 W=5.4e-07 AD=3.313e-13 AS=2.592e-13 PD=1.95333e-06 PS=2.04e-06 $X=1620 $Y=1480 $dt=0
M2 gnd3i! B 8 gnd3i! ne3i L=3.5e-07 W=5.4e-07 AD=2.92808e-13 AS=3.313e-13 PD=1.47273e-06 PS=1.95333e-06 $X=2450 $Y=1010 $dt=0
M3 Q 9 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=4.82592e-13 PD=2.74e-06 PS=2.42727e-06 $X=3510 $Y=660 $dt=0
M4 9 C vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=2.295e-13 AS=1.03315e-12 PD=1.39e-06 PS=4.25e-06 $X=975 $Y=2880 $dt=1
M5 10 A 9 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=2.295e-13 PD=1.1e-06 PS=1.39e-06 $X=1815 $Y=2880 $dt=1
M6 vdd3i! B 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.77448e-13 AS=1.0625e-13 PD=1.94425e-06 PS=1.1e-06 $X=2365 $Y=2880 $dt=1
M7 Q 9 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=7.92002e-13 PD=3.78e-06 PS=3.22516e-06 $X=3560 $Y=2410 $dt=1
.ends OA21JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: EO2JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt EO2JI3VX0 vdd3i! gnd3i! B A Q
*.DEVICECLIMB
** N=10 EP=5 FDC=10
M0 8 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.628e-13 PD=9.6e-07 PS=3.52e-06 $X=660 $Y=1130 $dt=0
M1 gnd3i! A 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.0445e-13 AS=1.134e-13 PD=1.34e-06 PS=9.6e-07 $X=1550 $Y=1130 $dt=0
M2 7 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.25e-14 AS=2.0445e-13 PD=6.7e-07 PS=1.34e-06 $X=2670 $Y=980 $dt=0
M3 Q A 7 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.503e-13 AS=5.25e-14 PD=1.15e-06 PS=6.7e-07 $X=3270 $Y=980 $dt=0
M4 gnd3i! 8 Q gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.0464e-12 AS=1.503e-13 PD=4.3e-06 PS=1.15e-06 $X=4200 $Y=1130 $dt=0
M5 10 B vdd3i! vdd3i! pe3i L=3e-07 W=9e-07 AD=1.35e-13 AS=7.175e-13 PD=1.2e-06 PS=4.61e-06 $X=575 $Y=2410 $dt=1
M6 8 A 10 vdd3i! pe3i L=3e-07 W=9e-07 AD=5.38188e-13 AS=1.35e-13 PD=3.13778e-06 PS=1.2e-06 $X=1175 $Y=2410 $dt=1
M7 vdd3i! B 9 vdd3i! pe3i L=3e-07 W=1.3e-06 AD=5.321e-13 AS=5.76588e-13 PD=2.43e-06 PS=3.57778e-06 $X=2795 $Y=2520 $dt=1
M8 9 A vdd3i! vdd3i! pe3i L=3e-07 W=1.3e-06 AD=3.835e-13 AS=5.321e-13 PD=1.89e-06 PS=2.43e-06 $X=3765 $Y=2410 $dt=1
M9 Q 8 9 vdd3i! pe3i L=3e-07 W=1.3e-06 AD=6.565e-13 AS=3.835e-13 PD=3.61e-06 PS=1.89e-06 $X=4655 $Y=2410 $dt=1
.ends EO2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO3JI3VX0                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO3JI3VX0 vdd3i! gnd3i! C Q B A
*.DEVICECLIMB
** N=9 EP=6 FDC=6
M0 Q C gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=5.75467e-13 PD=9.6e-07 PS=2.95333e-06 $X=615 $Y=1130 $dt=0
M1 gnd3i! B Q gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=5.75467e-13 AS=1.134e-13 PD=2.95333e-06 PS=9.6e-07 $X=1505 $Y=1130 $dt=0
M2 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=5.75467e-13 PD=1.8e-06 PS=2.95333e-06 $X=2390 $Y=1130 $dt=0
M3 9 C vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=1.55e-13 AS=1.3584e-12 PD=1.31e-06 PS=5.15e-06 $X=955 $Y=2410 $dt=1
M4 8 B 9 vdd3i! pe3i L=3e-07 W=1e-06 AD=1.55e-13 AS=1.55e-13 PD=1.31e-06 PS=1.31e-06 $X=1565 $Y=2410 $dt=1
M5 Q A 8 vdd3i! pe3i L=3e-07 W=1e-06 AD=4.8e-13 AS=1.55e-13 PD=2.96e-06 PS=1.31e-06 $X=2175 $Y=2410 $dt=1
.ends NO3JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AN31JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AN31JI3VX1 vdd3i! gnd3i! A B C Q D
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 10 A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.335e-13 AS=6.098e-13 PD=1.19e-06 PS=3.52e-06 $X=660 $Y=660 $dt=0
M1 9 B 10 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.35725e-13 AS=1.335e-13 PD=1.195e-06 PS=1.19e-06 $X=1310 $Y=660 $dt=0
M2 Q C 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.0257e-13 AS=1.35725e-13 PD=1.8043e-06 PS=1.195e-06 $X=1965 $Y=660 $dt=0
M3 gnd3i! D Q gnd3i! ne3i L=3.5e-07 W=5.75e-07 AD=5.783e-13 AS=1.9548e-13 PD=3.52e-06 PS=1.1657e-06 $X=2910 $Y=975 $dt=0
M4 11 A vdd3i! vdd3i! pe3i L=3.00061e-07 W=1.44471e-06 AD=3.0525e-13 AS=5.93475e-13 PD=1.86471e-06 PS=3.72971e-06 $X=525 $Y=2425 $dt=1
M5 vdd3i! B 11 vdd3i! pe3i L=3.00061e-07 W=1.44471e-06 AD=4.42387e-13 AS=3.0525e-13 PD=2.08971e-06 PS=1.86471e-06 $X=1365 $Y=2425 $dt=1
M6 11 C vdd3i! vdd3i! pe3i L=3.00061e-07 W=1.44471e-06 AD=2.6565e-13 AS=4.42387e-13 PD=1.86471e-06 PS=2.08971e-06 $X=2310 $Y=2425 $dt=1
M7 Q D 11 vdd3i! pe3i L=3.00061e-07 W=1.44471e-06 AD=7.2375e-13 AS=2.6565e-13 PD=3.85971e-06 PS=1.86471e-06 $X=2910 $Y=2425 $dt=1
.ends AN31JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND2JI3VX0                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND2JI3VX0 vdd3i! gnd3i! A B Q
*.DEVICECLIMB
** N=8 EP=5 FDC=6
M0 7 A 8 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=7e-14 AS=2.688e-13 PD=8.1e-07 PS=2.08e-06 $X=820 $Y=990 $dt=0
M1 gnd3i! B 7 gnd3i! ne3i L=3.5e-07 W=5.6e-07 AD=3.536e-13 AS=7e-14 PD=2.12571e-06 PS=8.1e-07 $X=1420 $Y=990 $dt=0
M2 Q 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=2.016e-13 AS=2.652e-13 PD=1.8e-06 PS=1.59429e-06 $X=2390 $Y=1130 $dt=0
M3 8 A vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=1.89e-13 AS=7.276e-13 PD=1.24e-06 PS=4.56e-06 $X=580 $Y=2410 $dt=1
M4 vdd3i! B 8 vdd3i! pe3i L=3e-07 W=7e-07 AD=5.276e-13 AS=1.89e-13 PD=2.48e-06 PS=1.24e-06 $X=1420 $Y=2410 $dt=1
M5 Q 8 vdd3i! vdd3i! pe3i L=3e-07 W=7e-07 AD=3.36e-13 AS=5.276e-13 PD=2.36e-06 PS=2.48e-06 $X=2440 $Y=2410 $dt=1
.ends AND2JI3VX0

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO3I1JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO3I1JI3VX1 vdd3i! gnd3i! AN Q B C
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 gnd3i! AN 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.99484e-13 AS=2.016e-13 PD=1.19267e-06 PS=1.8e-06 $X=620 $Y=1130 $dt=0
M1 Q 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=4.22716e-13 PD=1.43e-06 PS=2.52733e-06 $X=1550 $Y=660 $dt=0
M2 gnd3i! B Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=2440 $Y=660 $dt=0
M3 Q C gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.272e-13 AS=3.494e-13 PD=2.74e-06 PS=1.86e-06 $X=3410 $Y=660 $dt=0
M4 vdd3i! AN 8 vdd3i! pe3i L=3e-07 W=7e-07 AD=4.49443e-13 AS=3.36e-13 PD=1.73175e-06 PS=2.36e-06 $X=620 $Y=2415 $dt=1
M5 10 8 vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=9.05307e-13 PD=1.72e-06 PS=3.48825e-06 $X=1770 $Y=2410 $dt=1
M6 9 B 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.1855e-13 AS=2.1855e-13 PD=1.72e-06 PS=1.72e-06 $X=2380 $Y=2410 $dt=1
M7 Q C 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=2.1855e-13 PD=3.78e-06 PS=1.72e-06 $X=2990 $Y=2410 $dt=1
.ends NO3I1JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AN211JI3VX1                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AN211JI3VX1 vdd3i! gnd3i! B A Q C D
*.DEVICECLIMB
** N=11 EP=7 FDC=8
M0 9 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=6.47e-13 PD=1.14e-06 PS=3.58e-06 $X=690 $Y=660 $dt=0
M1 Q A 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.9785e-13 AS=1.1125e-13 PD=1.71704e-06 PS=1.14e-06 $X=1290 $Y=660 $dt=0
M2 gnd3i! C Q gnd3i! ne3i L=3.5e-07 W=6.65e-07 AD=5.036e-13 AS=2.2255e-13 PD=2.145e-06 PS=1.28296e-06 $X=2250 $Y=885 $dt=0
M3 Q D gnd3i! gnd3i! ne3i L=3.5e-07 W=6.65e-07 AD=3.22525e-13 AS=5.036e-13 PD=2.3e-06 PS=2.145e-06 $X=3505 $Y=885 $dt=0
M4 vdd3i! B 11 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.5825e-13 AS=6.768e-13 PD=2.06e-06 PS=3.78e-06 $X=620 $Y=2410 $dt=1
M5 11 A vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=4.1595e-13 AS=4.5825e-13 PD=2e-06 PS=2.06e-06 $X=1570 $Y=2410 $dt=1
M6 10 C 11 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=2.115e-13 AS=4.1595e-13 PD=1.71e-06 PS=2e-06 $X=2460 $Y=2410 $dt=1
M7 Q D 10 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=6.768e-13 AS=2.115e-13 PD=3.78e-06 PS=1.71e-06 $X=3060 $Y=2410 $dt=1
.ends AN211JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO22JI3VX1                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO22JI3VX1 vdd3i! gnd3i! B A Q C
*.DEVICECLIMB
** N=10 EP=6 FDC=8
M0 8 B gnd3i! gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=1.134e-13 AS=4.87734e-13 PD=9.6e-07 PS=2.24324e-06 $X=720 $Y=1130 $dt=0
M1 gnd3i! A 8 gnd3i! ne3i L=3.5e-07 W=4.2e-07 AD=4.87734e-13 AS=1.134e-13 PD=2.24324e-06 PS=9.6e-07 $X=1610 $Y=1130 $dt=0
M2 Q 8 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=1.03353e-12 PD=1.43e-06 PS=4.75353e-06 $X=2580 $Y=660 $dt=0
M3 gnd3i! C Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=6.098e-13 AS=2.403e-13 PD=3.52e-06 PS=1.43e-06 $X=3470 $Y=660 $dt=0
M4 10 B vdd3i! vdd3i! pe3i L=3e-07 W=8.5e-07 AD=1.0625e-13 AS=1.0178e-12 PD=1.1e-06 PS=4.78e-06 $X=770 $Y=2410 $dt=1
M5 8 A 10 vdd3i! pe3i L=3e-07 W=8.5e-07 AD=4.505e-13 AS=1.0625e-13 PD=2.76e-06 PS=1.1e-06 $X=1320 $Y=2410 $dt=1
M6 9 8 Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=6.768e-13 PD=1.66e-06 PS=3.78e-06 $X=2920 $Y=2410 $dt=1
M7 vdd3i! C 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=9.682e-13 AS=1.7625e-13 PD=4.66e-06 PS=1.66e-06 $X=3470 $Y=2410 $dt=1
.ends NO22JI3VX1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA2JI3VX2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA2JI3VX2 vdd3i! gnd3i! B Q A
*.DEVICECLIMB
** N=8 EP=5 FDC=8
M0 8 B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=7.09e-13 PD=1.14e-06 PS=3.68e-06 $X=740 $Y=660 $dt=0
M1 Q A 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=1.1125e-13 PD=1.43e-06 PS=1.14e-06 $X=1340 $Y=660 $dt=0
M2 7 A Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=2.403e-13 PD=1.14e-06 PS=1.43e-06 $X=2230 $Y=660 $dt=0
M3 gnd3i! B 7 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=7.09e-13 AS=1.1125e-13 PD=3.68e-06 PS=1.14e-06 $X=2830 $Y=660 $dt=0
M4 Q B vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.7e-13 AS=8.172e-13 PD=1.54e-06 PS=4.22e-06 $X=540 $Y=2410 $dt=1
M5 vdd3i! A Q vdd3i! pe3i L=3e-07 W=1e-06 AD=8.172e-13 AS=2.7e-13 PD=4.22e-06 PS=1.54e-06 $X=1380 $Y=2410 $dt=1
M6 Q A vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.7e-13 AS=8.172e-13 PD=1.54e-06 PS=4.22e-06 $X=2240 $Y=2410 $dt=1
M7 vdd3i! B Q vdd3i! pe3i L=3e-07 W=1e-06 AD=8.172e-13 AS=2.7e-13 PD=4.22e-06 PS=1.54e-06 $X=3080 $Y=2410 $dt=1
.ends NA2JI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NO2JI3VX2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NO2JI3VX2 vdd3i! gnd3i! B A Q
*.DEVICECLIMB
** N=8 EP=5 FDC=8
M0 Q B gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=6.842e-13 PD=1.43e-06 PS=3.64e-06 $X=720 $Y=660 $dt=0
M1 gnd3i! A Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=3.494e-13 AS=2.403e-13 PD=1.86e-06 PS=1.43e-06 $X=1610 $Y=660 $dt=0
M2 Q A gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.403e-13 AS=3.494e-13 PD=1.43e-06 PS=1.86e-06 $X=2580 $Y=660 $dt=0
M3 gnd3i! B Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=6.098e-13 AS=2.403e-13 PD=3.52e-06 PS=1.43e-06 $X=3470 $Y=660 $dt=0
M4 8 B vdd3i! vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=1.6898e-12 PD=1.66e-06 PS=5.48e-06 $X=1120 $Y=2410 $dt=1
M5 Q A 8 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=3.807e-13 AS=1.7625e-13 PD=1.95e-06 PS=1.66e-06 $X=1670 $Y=2410 $dt=1
M6 7 A Q vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.7625e-13 AS=3.807e-13 PD=1.66e-06 PS=1.95e-06 $X=2510 $Y=2410 $dt=1
M7 vdd3i! B 7 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=1.6898e-12 AS=1.7625e-13 PD=5.48e-06 PS=1.66e-06 $X=3060 $Y=2410 $dt=1
.ends NO2JI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NA2I1JI3VX2                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NA2I1JI3VX2 vdd3i! gnd3i! AN Q B
*.DEVICECLIMB
** N=9 EP=5 FDC=10
M0 gnd3i! AN 9 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=4.672e-13 AS=4.272e-13 PD=2.05e-06 PS=2.74e-06 $X=620 $Y=660 $dt=0
M1 8 9 gnd3i! gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=4.672e-13 PD=1.14e-06 PS=2.05e-06 $X=1780 $Y=660 $dt=0
M2 Q B 8 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=2.759e-13 AS=1.1125e-13 PD=1.51e-06 PS=1.14e-06 $X=2380 $Y=660 $dt=0
M3 7 B Q gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=1.1125e-13 AS=2.759e-13 PD=1.14e-06 PS=1.51e-06 $X=3350 $Y=660 $dt=0
M4 gnd3i! 9 7 gnd3i! ne3i L=3.5e-07 W=8.9e-07 AD=7.09e-13 AS=1.1125e-13 PD=3.68e-06 PS=1.14e-06 $X=3950 $Y=660 $dt=0
M5 vdd3i! AN 9 vdd3i! pe3i L=3e-07 W=1.41e-06 AD=9.9878e-13 AS=6.768e-13 PD=4.57664e-06 PS=3.78e-06 $X=620 $Y=2410 $dt=1
M6 Q 9 vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.7e-13 AS=7.08355e-13 PD=1.54e-06 PS=3.24584e-06 $X=1540 $Y=2410 $dt=1
M7 vdd3i! B Q vdd3i! pe3i L=3e-07 W=1e-06 AD=7.08355e-13 AS=2.7e-13 PD=3.24584e-06 PS=1.54e-06 $X=2380 $Y=2410 $dt=1
M8 Q B vdd3i! vdd3i! pe3i L=3e-07 W=1e-06 AD=2.7e-13 AS=7.08355e-13 PD=1.54e-06 PS=3.24584e-06 $X=3280 $Y=2410 $dt=1
M9 vdd3i! 9 Q vdd3i! pe3i L=3e-07 W=1e-06 AD=7.08355e-13 AS=2.7e-13 PD=3.24584e-06 PS=1.54e-06 $X=4120 $Y=2410 $dt=1
.ends NA2I1JI3VX2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP25JI3V                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP25JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=12
M0 gnd3i! 5 4 gnd3i! ne3i L=3.5e-07 W=8.8e-07 AD=2.376e-13 AS=4.224e-13 PD=1.42e-06 PS=2.72e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=1510 $Y=660 $dt=0
M2 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=3990 $Y=660 $dt=0
M3 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=6470 $Y=660 $dt=0
M4 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=8950 $Y=660 $dt=0
M5 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.94e-06 W=8.8e-07 AD=4.312e-13 AS=2.376e-13 PD=2.74e-06 PS=1.42e-06 $X=11430 $Y=660 $dt=0
M6 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.5505e-13 AS=6.312e-13 PD=1.855e-06 PS=3.59e-06 $X=620 $Y=2505 $dt=1
M7 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.5505e-13 AS=3.5505e-13 PD=1.855e-06 PS=1.855e-06 $X=3090 $Y=2505 $dt=1
M8 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.5505e-13 AS=3.5505e-13 PD=1.855e-06 PS=1.855e-06 $X=5560 $Y=2505 $dt=1
M9 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.5505e-13 AS=3.5505e-13 PD=1.855e-06 PS=1.855e-06 $X=8030 $Y=2505 $dt=1
M10 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.93e-06 W=1.315e-06 AD=3.84638e-13 AS=3.5505e-13 PD=1.9e-06 PS=1.855e-06 $X=10500 $Y=2505 $dt=1
M11 5 4 vdd3i! vdd3i! pe3i L=3e-07 W=1.315e-06 AD=7.56575e-13 AS=3.84638e-13 PD=3.91e-06 PS=1.9e-06 $X=13015 $Y=2505 $dt=1
.ends DECAP25JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP10JI3V                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP10JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=6
M0 gnd3i! 5 4 gnd3i! ne3i L=3.5e-07 W=8.8e-07 AD=2.376e-13 AS=4.224e-13 PD=1.42e-06 PS=2.72e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.445e-06 W=8.8e-07 AD=2.376e-13 AS=2.376e-13 PD=1.42e-06 PS=1.42e-06 $X=1510 $Y=660 $dt=0
M2 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.445e-06 W=8.8e-07 AD=6.046e-13 AS=2.376e-13 PD=3.5e-06 PS=1.42e-06 $X=3495 $Y=660 $dt=0
M3 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.425e-06 W=1.315e-06 AD=3.5505e-13 AS=8.308e-13 PD=1.855e-06 PS=4.37e-06 $X=660 $Y=2505 $dt=1
M4 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.425e-06 W=1.315e-06 AD=3.71488e-13 AS=3.5505e-13 PD=1.88e-06 PS=1.855e-06 $X=2625 $Y=2505 $dt=1
M5 5 4 vdd3i! vdd3i! pe3i L=3e-07 W=1.315e-06 AD=7.56575e-13 AS=3.71488e-13 PD=3.91e-06 PS=1.88e-06 $X=4615 $Y=2505 $dt=1
.ends DECAP10JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP7JI3V                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP7JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=4
M0 gnd3i! 5 4 gnd3i! ne3i L=3.5e-07 W=8.8e-07 AD=2.376e-13 AS=4.224e-13 PD=1.42e-06 PS=2.72e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.75e-06 W=8.8e-07 AD=6.046e-13 AS=2.376e-13 PD=3.5e-06 PS=1.42e-06 $X=1510 $Y=660 $dt=0
M2 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.71e-06 W=1.315e-06 AD=3.87925e-13 AS=8.308e-13 PD=1.905e-06 PS=4.37e-06 $X=660 $Y=2505 $dt=1
M3 5 4 vdd3i! vdd3i! pe3i L=3e-07 W=1.315e-06 AD=7.237e-13 AS=3.87925e-13 PD=3.86e-06 PS=1.905e-06 $X=2960 $Y=2505 $dt=1
.ends DECAP7JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP5JI3V                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP5JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=2
M0 gnd3i! 5 4 gnd3i! ne3i L=1.48e-06 W=8.3e-07 AD=5.786e-13 AS=4.568e-13 PD=3.4e-06 PS=2.82e-06 $X=660 $Y=660 $dt=0
M1 5 4 vdd3i! vdd3i! pe3i L=1.46e-06 W=1.36e-06 AD=7.564e-13 AS=8.542e-13 PD=3.9e-06 PS=4.46e-06 $X=660 $Y=2460 $dt=1
.ends DECAP5JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: DECAP15JI3V                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt DECAP15JI3V vdd3i! gnd3i!
*.DEVICECLIMB
** N=5 EP=2 FDC=8
M0 gnd3i! 5 4 gnd3i! ne3i L=3.5e-07 W=8.8e-07 AD=2.42e-13 AS=4.224e-13 PD=1.43e-06 PS=2.72e-06 $X=620 $Y=660 $dt=0
M1 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.71e-06 W=8.8e-07 AD=2.42e-13 AS=2.42e-13 PD=1.43e-06 PS=1.43e-06 $X=1520 $Y=660 $dt=0
M2 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.71e-06 W=8.8e-07 AD=2.376e-13 AS=2.42e-13 PD=1.42e-06 PS=1.43e-06 $X=3780 $Y=660 $dt=0
M3 gnd3i! 5 gnd3i! gnd3i! ne3i L=1.71e-06 W=8.8e-07 AD=6.046e-13 AS=2.376e-13 PD=3.5e-06 PS=1.42e-06 $X=6030 $Y=660 $dt=0
M4 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.7e-06 W=1.315e-06 AD=3.5505e-13 AS=8.308e-13 PD=1.855e-06 PS=4.37e-06 $X=660 $Y=2505 $dt=1
M5 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.7e-06 W=1.315e-06 AD=3.5505e-13 AS=3.5505e-13 PD=1.855e-06 PS=1.855e-06 $X=2900 $Y=2505 $dt=1
M6 vdd3i! 4 vdd3i! vdd3i! pe3i L=1.7e-06 W=1.315e-06 AD=3.78063e-13 AS=3.5505e-13 PD=1.89e-06 PS=1.855e-06 $X=5140 $Y=2505 $dt=1
M7 5 4 vdd3i! vdd3i! pe3i L=3e-07 W=1.315e-06 AD=7.56575e-13 AS=3.78063e-13 PD=3.91e-06 PS=1.89e-06 $X=7415 $Y=2505 $dt=1
.ends DECAP15JI3V

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: aska_dig                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt aska_dig DAC<0> DAC<1> DAC<2> DAC<3> DAC<4> DAC<5> IC_addr<0> IC_addr<1> SPI_CS SPI_Clk
+ SPI_MOSI clk down_switches<0> down_switches<10> down_switches<11> down_switches<12> down_switches<13> down_switches<14> down_switches<15> down_switches<16>
+ down_switches<17> down_switches<18> down_switches<19> down_switches<1> down_switches<20> down_switches<21> down_switches<22> down_switches<23> down_switches<24> down_switches<25>
+ down_switches<26> down_switches<27> down_switches<28> down_switches<29> down_switches<2> down_switches<30> down_switches<31> down_switches<3> down_switches<4> down_switches<5>
+ down_switches<6> down_switches<7> down_switches<8> down_switches<9> enable porborn pulse_active reset_l up_switches<0> up_switches<10>
+ up_switches<11> up_switches<12> up_switches<13> up_switches<14> up_switches<15> up_switches<16> up_switches<17> up_switches<18> up_switches<19> up_switches<1>
+ up_switches<20> up_switches<21> up_switches<22> up_switches<23> up_switches<24> up_switches<25> up_switches<26> up_switches<27> up_switches<28> up_switches<29>
+ up_switches<2> up_switches<30> up_switches<31> up_switches<3> up_switches<4> up_switches<5> up_switches<6> up_switches<7> up_switches<8> up_switches<9>
** N=1450 EP=80 FDC=26859
X8323 3 1 69 66 BUJI3VX2 $T=174160 87360 1 0 $X=173730 $Y=82240
X8324 3 1 570 up_switches<31> BUJI3VX2 $T=246960 24640 0 180 $X=243170 $Y=19520
X8325 3 1 1102 up_switches<30> BUJI3VX2 $T=250320 24640 0 180 $X=246530 $Y=19520
X8326 3 1 1249 up_switches<29> BUJI3VX2 $T=250880 24640 1 0 $X=250450 $Y=19520
X8327 3 1 578 518 BUJI3VX2 $T=252560 159040 0 0 $X=252130 $Y=158400
X8328 3 1 966 up_switches<28> BUJI3VX2 $T=254240 24640 1 0 $X=253810 $Y=19520
X8329 3 1 607 536 BUJI3VX2 $T=256480 203840 0 0 $X=256050 $Y=203200
X8330 3 1 104 up_switches<27> BUJI3VX2 $T=257600 24640 1 0 $X=257170 $Y=19520
X8331 3 1 571 up_switches<26> BUJI3VX2 $T=260960 24640 1 0 $X=260530 $Y=19520
X8332 3 1 575 up_switches<25> BUJI3VX2 $T=264880 24640 1 0 $X=264450 $Y=19520
X8333 3 1 107 130 BUJI3VX2 $T=266000 33600 0 0 $X=265570 $Y=32960
X8334 3 1 567 up_switches<24> BUJI3VX2 $T=268240 24640 1 0 $X=267810 $Y=19520
X8335 3 1 clk 12 BUJI3VX2 $T=273280 212800 0 180 $X=269490 $Y=207680
X8336 3 1 578 131 BUJI3VX2 $T=273840 185920 1 0 $X=273410 $Y=180800
X8337 3 1 904 up_switches<23> BUJI3VX2 $T=277760 24640 1 0 $X=277330 $Y=19520
X8338 3 1 589 up_switches<21> BUJI3VX2 $T=285040 24640 1 0 $X=284610 $Y=19520
X8339 3 1 612 up_switches<20> BUJI3VX2 $T=288960 24640 1 0 $X=288530 $Y=19520
X8340 3 1 602 up_switches<19> BUJI3VX2 $T=292320 24640 1 0 $X=291890 $Y=19520
X8341 3 1 1263 643 BUJI3VX2 $T=299040 212800 0 0 $X=298610 $Y=212160
X8342 3 1 131 154 BUJI3VX2 $T=371840 123200 0 0 $X=371410 $Y=122560
X8343 3 1 668 1010 1008 AND2JI3VX1 $T=67200 24640 1 180 $X=63410 $Y=24000
X8344 3 1 668 1215 1381 AND2JI3VX1 $T=68880 24640 0 0 $X=68450 $Y=24000
X8345 3 1 668 253 1016 AND2JI3VX1 $T=76720 33600 0 180 $X=72930 $Y=28480
X8346 3 1 668 257 1029 AND2JI3VX1 $T=84000 33600 0 180 $X=80210 $Y=28480
X8347 3 1 668 276 1033 AND2JI3VX1 $T=89040 33600 0 180 $X=85250 $Y=28480
X8348 3 1 668 822 1043 AND2JI3VX1 $T=93520 24640 0 0 $X=93090 $Y=24000
X8349 3 1 242 208 790 EN2JI3VX0 $T=70000 176960 1 180 $X=63970 $Y=176320
X8350 3 1 265 1031 1028 EN2JI3VX0 $T=84560 203840 0 180 $X=78530 $Y=198720
X8351 3 1 274 282 814 EN2JI3VX0 $T=91280 194880 1 180 $X=85250 $Y=194240
X8352 3 1 965 474 1238 EN2JI3VX0 $T=204400 194880 0 180 $X=198370 $Y=189760
X8353 3 1 1084 484 1088 EN2JI3VX0 $T=205520 212800 1 0 $X=205090 $Y=207680
X8354 3 1 603 1117 1382 EN2JI3VX0 $T=276640 221760 0 180 $X=270610 $Y=216640
X8355 3 1 935 937 934 EN2JI3VX0 $T=343280 203840 0 180 $X=337250 $Y=198720
X8356 3 1 958 1383 1297 NA2I1JI3VX1 $T=53760 203840 1 0 $X=53330 $Y=198720
X8357 3 1 1003 1005 221 NA2I1JI3VX1 $T=58800 185920 0 0 $X=58370 $Y=185280
X8358 3 1 228 221 794 NA2I1JI3VX1 $T=62160 185920 0 0 $X=61730 $Y=185280
X8359 3 1 227 22 278 NA2I1JI3VX1 $T=64960 203840 1 0 $X=64530 $Y=198720
X8360 3 1 794 212 228 NA2I1JI3VX1 $T=68880 185920 1 180 $X=65090 $Y=185280
X8361 3 1 1019 1024 1017 NA2I1JI3VX1 $T=72800 105280 1 0 $X=72370 $Y=100160
X8362 3 1 323 1017 256 NA2I1JI3VX1 $T=79520 105280 0 180 $X=75730 $Y=100160
X8363 3 1 1020 277 807 NA2I1JI3VX1 $T=77280 185920 1 0 $X=76850 $Y=180800
X8364 3 1 1015 272 265 NA2I1JI3VX1 $T=78400 194880 1 0 $X=77970 $Y=189760
X8365 3 1 265 807 1015 NA2I1JI3VX1 $T=85120 194880 0 180 $X=81330 $Y=189760
X8366 3 1 1031 281 265 NA2I1JI3VX1 $T=83440 203840 0 0 $X=83010 $Y=203200
X8367 3 1 33 1042 270 NA2I1JI3VX1 $T=94080 105280 1 180 $X=90290 $Y=104640
X8368 3 1 278 813 1041 NA2I1JI3VX1 $T=91840 203840 1 0 $X=91410 $Y=198720
X8369 3 1 824 823 49 NA2I1JI3VX1 $T=96880 185920 1 0 $X=96450 $Y=180800
X8370 3 1 296 825 1042 NA2I1JI3VX1 $T=101920 105280 1 180 $X=98130 $Y=104640
X8371 3 1 829 35 294 NA2I1JI3VX1 $T=104720 194880 0 180 $X=100930 $Y=189760
X8372 3 1 348 346 834 NA2I1JI3VX1 $T=135520 185920 1 180 $X=131730 $Y=185280
X8373 3 1 847 1058 853 NA2I1JI3VX1 $T=148960 203840 1 0 $X=148530 $Y=198720
X8374 3 1 1344 1345 416 NA2I1JI3VX1 $T=166320 203840 0 180 $X=162530 $Y=198720
X8375 3 1 484 498 1084 NA2I1JI3VX1 $T=204400 194880 0 0 $X=203970 $Y=194240
X8376 3 1 498 100 885 NA2I1JI3VX1 $T=219520 194880 1 0 $X=219090 $Y=189760
X8377 3 1 98 493 885 NA2I1JI3VX1 $T=225680 185920 1 180 $X=221890 $Y=185280
X8378 3 1 516 1093 97 NA2I1JI3VX1 $T=232400 185920 0 180 $X=228610 $Y=180800
X8379 3 1 1133 923 142 NA2I1JI3VX1 $T=313040 168000 0 0 $X=312610 $Y=167360
X8380 3 1 142 697 1133 NA2I1JI3VX1 $T=328720 168000 1 180 $X=324930 $Y=167360
X8381 3 1 926 698 142 NA2I1JI3VX1 $T=325360 194880 1 0 $X=324930 $Y=189760
X8382 3 1 937 1141 935 NA2I1JI3VX1 $T=337120 194880 0 180 $X=333330 $Y=189760
X8383 3 1 942 940 727 NA2I1JI3VX1 $T=343280 194880 1 0 $X=342850 $Y=189760
X8384 3 1 252 246 805 24 NO3I2JI3VX1 $T=78400 194880 1 180 $X=74050 $Y=194240
X8385 3 1 292 246 46 235 NO3I2JI3VX1 $T=100240 194880 0 180 $X=95890 $Y=189760
X8386 3 1 313 enable 314 1221 NO3I2JI3VX1 $T=117040 185920 0 180 $X=112690 $Y=180800
X8387 3 1 1050 246 314 368 NO3I2JI3VX1 $T=126000 194880 1 0 $X=125570 $Y=189760
X8388 3 1 1238 493 1313 1384 NO3I2JI3VX1 $T=203280 185920 1 180 $X=198930 $Y=185280
X8389 3 1 1134 936 729 929 NO3I2JI3VX1 $T=327040 176960 1 0 $X=326610 $Y=171840
X8390 3 1 reset_l 488 494 NA2JI3VX1 $T=208320 221760 1 0 $X=207890 $Y=216640
X8391 3 1 12 69 BUJI3VX1 $T=52640 24640 0 0 $X=52210 $Y=24000
X8392 3 1 661 514 BUJI3VX1 $T=66640 141120 0 0 $X=66210 $Y=140480
X8393 3 1 55 490 BUJI3VX1 $T=207200 42560 1 0 $X=206770 $Y=37440
X8394 3 1 514 891 BUJI3VX1 $T=230160 69440 0 0 $X=229730 $Y=68800
X8395 3 1 SPI_Clk 661 BUJI3VX1 $T=309120 105280 0 0 $X=308690 $Y=104640
X8396 3 1 180 974 14 191 DFRRQJI3VX4 $T=23520 60480 1 0 $X=23090 $Y=55360
X8397 3 1 180 789 14 244 DFRRQJI3VX4 $T=59920 42560 1 0 $X=59490 $Y=37440
X8398 3 1 180 1030 14 276 DFRRQJI3VX4 $T=76720 87360 0 0 $X=76290 $Y=86720
X8399 3 1 185 1051 4 348 DFRRQJI3VX4 $T=122640 212800 1 0 $X=122210 $Y=207680
X8400 3 1 618 635 116 620 DFRRQJI3VX4 $T=302400 221760 0 180 $X=284050 $Y=216640
X8401 3 1 161 1275 111 687 DFRRQJI3VX4 $T=344400 212800 1 180 $X=326050 $Y=212160
X8402 3 1 161 1276 111 701 DFRRQJI3VX4 $T=344960 212800 0 180 $X=326610 $Y=207680
X8403 3 1 161 715 111 935 DFRRQJI3VX4 $T=355040 203840 1 180 $X=336690 $Y=203200
X8404 3 1 161 743 111 945 DFRRQJI3VX4 $T=374080 185920 0 180 $X=355730 $Y=180800
X8405 3 1 1204 1332 BUJI3VX0 $T=30240 33600 1 0 $X=29810 $Y=28480
X8406 3 1 184 1334 BUJI3VX0 $T=34160 168000 0 0 $X=33730 $Y=167360
X8407 3 1 227 1385 BUJI3VX0 $T=38640 203840 1 0 $X=38210 $Y=198720
X8408 3 1 10 193 BUJI3VX0 $T=40320 33600 0 0 $X=39890 $Y=32960
X8409 3 1 201 773 BUJI3VX0 $T=50960 168000 1 0 $X=50530 $Y=162880
X8410 3 1 199 1207 BUJI3VX0 $T=52080 203840 0 0 $X=51650 $Y=203200
X8411 3 1 257 1217 BUJI3VX0 $T=75040 96320 1 0 $X=74610 $Y=91200
X8412 3 1 1041 269 BUJI3VX0 $T=86800 203840 0 0 $X=86370 $Y=203200
X8413 3 1 822 1219 BUJI3VX0 $T=92400 96320 0 0 $X=91970 $Y=95680
X8414 3 1 369 839 BUJI3VX0 $T=140560 212800 1 0 $X=140130 $Y=207680
X8415 3 1 426 416 BUJI3VX0 $T=146160 203840 1 0 $X=145730 $Y=198720
X8416 3 1 852 853 BUJI3VX0 $T=150640 203840 0 0 $X=150210 $Y=203200
X8417 3 1 442 863 BUJI3VX0 $T=169680 221760 1 0 $X=169250 $Y=216640
X8418 3 1 597 322 BUJI3VX0 $T=185920 132160 0 180 $X=182690 $Y=127040
X8419 3 1 488 80 BUJI3VX0 $T=197120 212800 0 0 $X=196690 $Y=212160
X8420 3 1 porborn 480 BUJI3VX0 $T=205520 221760 1 0 $X=205090 $Y=216640
X8421 3 1 SPI_CS 565 BUJI3VX0 $T=218960 221760 1 0 $X=218530 $Y=216640
X8422 3 1 542 1315 BUJI3VX0 $T=243040 212800 0 0 $X=242610 $Y=212160
X8423 3 1 80 113 BUJI3VX0 $T=245840 212800 0 0 $X=245410 $Y=212160
X8424 3 1 SPI_MOSI 551 BUJI3VX0 $T=247520 221760 1 0 $X=247090 $Y=216640
X8425 3 1 648 503 BUJI3VX0 $T=250320 221760 1 0 $X=249890 $Y=216640
X8426 3 1 522 533 BUJI3VX0 $T=252000 194880 1 0 $X=251570 $Y=189760
X8427 3 1 559 562 BUJI3VX0 $T=253680 203840 0 0 $X=253250 $Y=203200
X8428 3 1 1114 1250 BUJI3VX0 $T=254800 168000 0 0 $X=254370 $Y=167360
X8429 3 1 598 900 BUJI3VX0 $T=255920 185920 1 0 $X=255490 $Y=180800
X8430 3 1 536 578 BUJI3VX0 $T=262640 176960 0 0 $X=262210 $Y=176320
X8431 3 1 536 108 BUJI3VX0 $T=263200 203840 0 0 $X=262770 $Y=203200
X8432 3 1 1382 1254 BUJI3VX0 $T=268240 221760 1 0 $X=267810 $Y=216640
X8433 3 1 580 1319 BUJI3VX0 $T=273280 185920 0 0 $X=272850 $Y=185280
X8434 3 1 119 1256 BUJI3VX0 $T=274400 176960 0 0 $X=273970 $Y=176320
X8435 3 1 597 172 BUJI3VX0 $T=277760 168000 1 0 $X=277330 $Y=162880
X8436 3 1 600 631 BUJI3VX0 $T=278320 221760 1 0 $X=277890 $Y=216640
X8437 3 1 1118 906 BUJI3VX0 $T=279440 194880 1 0 $X=279010 $Y=189760
X8438 3 1 643 607 BUJI3VX0 $T=281120 212800 0 0 $X=280690 $Y=212160
X8439 3 1 617 1120 BUJI3VX0 $T=285600 212800 1 0 $X=285170 $Y=207680
X8440 3 1 631 1263 BUJI3VX0 $T=294000 212800 1 0 $X=293570 $Y=207680
X8441 3 1 912 642 BUJI3VX0 $T=298480 194880 1 0 $X=298050 $Y=189760
X8442 3 1 1153 1283 BUJI3VX0 $T=349440 203840 1 0 $X=349010 $Y=198720
X8443 3 1 199 767 1386 227 AN21JI3VX1 $T=45360 203840 1 180 $X=41570 $Y=203200
X8444 3 1 107 768 6 196 AN21JI3VX1 $T=47040 69440 1 180 $X=43250 $Y=68800
X8445 3 1 239 783 1210 1161 AN21JI3VX1 $T=58800 194880 0 180 $X=55010 $Y=189760
X8446 3 1 55 778 213 18 AN21JI3VX1 $T=56560 42560 0 0 $X=56130 $Y=41920
X8447 3 1 22 786 252 1009 AN21JI3VX1 $T=60480 194880 0 0 $X=60050 $Y=194240
X8448 3 1 1017 29 1336 1019 AN21JI3VX1 $T=72800 105280 0 180 $X=69010 $Y=100160
X8449 3 1 282 36 820 819 AN21JI3VX1 $T=95760 185920 1 180 $X=91970 $Y=185280
X8450 3 1 1045 1042 283 296 AN21JI3VX1 $T=97440 105280 1 180 $X=93650 $Y=104640
X8451 3 1 282 1220 1387 1041 AN21JI3VX1 $T=95200 212800 0 0 $X=94770 $Y=212160
X8452 3 1 346 361 1050 54 AN21JI3VX1 $T=133280 194880 0 180 $X=129490 $Y=189760
X8453 3 1 369 353 1388 348 AN21JI3VX1 $T=136640 203840 1 180 $X=132850 $Y=203200
X8454 3 1 1304 387 1057 851 AN21JI3VX1 $T=155680 185920 0 180 $X=151890 $Y=180800
X8455 3 1 1229 368 847 362 AN21JI3VX1 $T=156800 203840 0 180 $X=153010 $Y=198720
X8456 3 1 63 368 1344 362 AN21JI3VX1 $T=162960 203840 0 180 $X=159170 $Y=198720
X8457 3 1 477 1311 1389 1313 AN21JI3VX1 $T=204400 185920 0 0 $X=203970 $Y=185280
X8458 3 1 97 1351 1390 1239 AN21JI3VX1 $T=222880 194880 1 0 $X=222450 $Y=189760
X8459 3 1 1352 86 890 508 AN21JI3VX1 $T=225680 203840 1 0 $X=225250 $Y=198720
X8460 3 1 894 895 1244 1372 AN21JI3VX1 $T=240800 185920 1 180 $X=237010 $Y=185280
X8461 3 1 701 1361 1270 687 AN21JI3VX1 $T=330960 203840 0 180 $X=327170 $Y=198720
X8462 3 1 155 690 1143 1144 AN21JI3VX1 $T=330960 185920 0 0 $X=330530 $Y=185280
X8463 3 1 1136 933 672 689 AN21JI3VX1 $T=335440 176960 1 0 $X=335010 $Y=171840
X8464 3 1 162 941 1391 939 AN21JI3VX1 $T=345520 176960 0 180 $X=341730 $Y=171840
X8465 3 1 225 8 996 1392 EN3JI3VX1 $T=43680 96320 1 0 $X=43250 $Y=91200
X8466 3 1 1005 1161 212 1393 NA3I2JI3VX1 $T=59360 194880 1 0 $X=58930 $Y=189760
X8467 3 1 1383 1009 22 1213 NA3I2JI3VX1 $T=60480 203840 1 0 $X=60050 $Y=198720
X8468 3 1 464 460 517 94 NA3I2JI3VX1 $T=188720 194880 0 0 $X=188290 $Y=194240
X8469 3 1 1093 1239 1353 1394 NA3I2JI3VX1 $T=227360 185920 0 0 $X=226930 $Y=185280
X8470 3 1 1395 1118 603 593 NA3I2JI3VX1 $T=277760 212800 0 180 $X=273410 $Y=207680
X8471 3 1 221 999 212 783 NA22JI3VX1 $T=54320 185920 0 0 $X=53890 $Y=185280
X8472 3 1 778 55 785 797 NA22JI3VX1 $T=61040 42560 0 0 $X=60610 $Y=41920
X8473 3 1 281 235 961 1038 NA22JI3VX1 $T=89600 203840 0 0 $X=89170 $Y=203200
X8474 3 1 383 1375 1168 361 NA22JI3VX1 $T=145600 194880 0 180 $X=141250 $Y=189760
X8475 3 1 840 846 377 403 NA22JI3VX1 $T=142240 185920 0 0 $X=141810 $Y=185280
X8476 3 1 863 362 861 445 NA22JI3VX1 $T=170800 203840 1 180 $X=166450 $Y=203200
X8477 3 1 498 86 489 508 NA22JI3VX1 $T=207760 194880 0 0 $X=207330 $Y=194240
X8478 3 1 926 672 enable 968 NA22JI3VX1 $T=313600 194880 0 0 $X=313170 $Y=194240
X8479 3 1 152 688 682 153 NA22JI3VX1 $T=333200 176960 1 180 $X=328850 $Y=176320
X8480 3 1 672 1141 enable 1272 NA22JI3VX1 $T=334880 194880 1 180 $X=330530 $Y=194240
X8481 3 1 942 672 enable 1279 NA22JI3VX1 $T=344960 194880 1 180 $X=340610 $Y=194240
X8482 3 1 1154 1330 167 718 NA22JI3VX1 $T=356160 176960 0 180 $X=351810 $Y=171840
X8483 3 1 217 771 203 774 16 AN22JI3VX1 $T=47040 51520 1 0 $X=46610 $Y=46400
X8484 3 1 1211 203 778 13 202 AN22JI3VX1 $T=56000 51520 0 180 $X=51650 $Y=46400
X8485 3 1 225 260 780 266 11 AN22JI3VX1 $T=64960 96320 1 180 $X=60610 $Y=95680
X8486 3 1 280 260 1006 266 782 AN22JI3VX1 $T=64960 105280 1 180 $X=60610 $Y=104640
X8487 3 1 215 260 791 266 20 AN22JI3VX1 $T=70000 96320 1 180 $X=65650 $Y=95680
X8488 3 1 794 1013 259 796 236 AN22JI3VX1 $T=67200 185920 1 0 $X=66770 $Y=180800
X8489 3 1 1035 34 1396 260 323 AN22JI3VX1 $T=85120 96320 1 180 $X=80770 $Y=95680
X8490 3 1 960 34 809 260 33 AN22JI3VX1 $T=90160 96320 1 180 $X=85810 $Y=95680
X8491 3 1 818 260 816 34 1302 AN22JI3VX1 $T=91280 105280 0 180 $X=86930 $Y=100160
X8492 3 1 451 292 961 46 enable AN22JI3VX1 $T=100240 194880 1 180 $X=95890 $Y=194240
X8493 3 1 846 388 848 394 395 AN22JI3VX1 $T=144480 194880 0 0 $X=144050 $Y=194240
X8494 3 1 374 76 609 107 389 AN22JI3VX1 $T=145040 24640 0 0 $X=144610 $Y=24000
X8495 3 1 1064 59 855 856 420 AN22JI3VX1 $T=160720 194880 1 180 $X=156370 $Y=194240
X8496 3 1 439 1075 424 448 1074 AN22JI3VX1 $T=176400 194880 0 180 $X=172050 $Y=189760
X8497 3 1 442 452 963 448 75 AN22JI3VX1 $T=179760 203840 1 0 $X=179330 $Y=198720
X8498 3 1 451 517 489 460 enable AN22JI3VX1 $T=184240 194880 0 0 $X=183810 $Y=194240
X8499 3 1 1244 1177 517 892 549 AN22JI3VX1 $T=236320 194880 0 180 $X=231970 $Y=189760
X8500 3 1 1258 649 746 130 910 AN22JI3VX1 $T=288400 33600 1 0 $X=287970 $Y=28480
X8501 3 1 629 649 740 130 1121 AN22JI3VX1 $T=295120 42560 0 180 $X=290770 $Y=37440
X8502 3 1 916 134 676 658 1128 AN22JI3VX1 $T=306320 168000 1 180 $X=301970 $Y=167360
X8503 3 1 1125 667 920 134 662 AN22JI3VX1 $T=304640 185920 0 0 $X=304210 $Y=185280
X8504 3 1 811 1298 DLY1JI3VX1 $T=53200 176960 1 0 $X=52770 $Y=171840
X8505 3 1 1209 214 DLY1JI3VX1 $T=53760 87360 0 0 $X=53330 $Y=86720
X8506 3 1 224 220 DLY1JI3VX1 $T=56560 69440 1 0 $X=56130 $Y=64320
X8507 3 1 230 223 DLY1JI3VX1 $T=58800 176960 1 0 $X=58370 $Y=171840
X8508 3 1 241 245 DLY1JI3VX1 $T=71120 42560 0 0 $X=70690 $Y=41920
X8509 3 1 427 804 DLY1JI3VX1 $T=73920 159040 0 0 $X=73490 $Y=158400
X8510 3 1 248 258 DLY1JI3VX1 $T=76720 51520 0 0 $X=76290 $Y=50880
X8511 3 1 1034 264 DLY1JI3VX1 $T=79520 159040 0 0 $X=79090 $Y=158400
X8512 3 1 262 267 DLY1JI3VX1 $T=82880 33600 0 0 $X=82450 $Y=32960
X8513 3 1 810 271 DLY1JI3VX1 $T=84000 176960 0 0 $X=83570 $Y=176320
X8514 3 1 324 305 DLY1JI3VX1 $T=88480 33600 0 0 $X=88050 $Y=32960
X8515 3 1 293 1367 DLY1JI3VX1 $T=89600 176960 0 0 $X=89170 $Y=176320
X8516 3 1 328 1039 DLY1JI3VX1 $T=99680 42560 1 180 $X=93650 $Y=41920
X8517 3 1 1044 1338 DLY1JI3VX1 $T=96880 24640 0 0 $X=96450 $Y=24000
X8518 3 1 301 300 DLY1JI3VX1 $T=105280 42560 1 180 $X=99250 $Y=41920
X8519 3 1 330 302 DLY1JI3VX1 $T=105280 87360 0 180 $X=99250 $Y=82240
X8520 3 1 371 827 DLY1JI3VX1 $T=105280 105280 0 180 $X=99250 $Y=100160
X8521 3 1 321 39 DLY1JI3VX1 $T=105280 150080 0 180 $X=99250 $Y=144960
X8522 3 1 325 42 DLY1JI3VX1 $T=113120 78400 1 0 $X=112690 $Y=73280
X8523 3 1 329 309 DLY1JI3VX1 $T=113120 78400 0 0 $X=112690 $Y=77760
X8524 3 1 366 310 DLY1JI3VX1 $T=113120 96320 0 0 $X=112690 $Y=95680
X8525 3 1 318 47 DLY1JI3VX1 $T=113120 150080 0 0 $X=112690 $Y=149440
X8526 3 1 327 315 DLY1JI3VX1 $T=116480 24640 0 0 $X=116050 $Y=24000
X8527 3 1 443 317 DLY1JI3VX1 $T=117600 123200 1 0 $X=117170 $Y=118080
X8528 3 1 831 832 DLY1JI3VX1 $T=118720 96320 0 0 $X=118290 $Y=95680
X8529 3 1 465 334 DLY1JI3VX1 $T=123200 123200 1 0 $X=122770 $Y=118080
X8530 3 1 51 335 DLY1JI3VX1 $T=123200 176960 0 0 $X=122770 $Y=176320
X8531 3 1 347 356 DLY1JI3VX1 $T=133840 33600 0 0 $X=133410 $Y=32960
X8532 3 1 381 357 DLY1JI3VX1 $T=133840 69440 0 0 $X=133410 $Y=68800
X8533 3 1 440 365 DLY1JI3VX1 $T=137760 114240 0 0 $X=137330 $Y=113600
X8534 3 1 472 367 DLY1JI3VX1 $T=138320 132160 0 0 $X=137890 $Y=131520
X8535 3 1 446 382 DLY1JI3VX1 $T=142800 141120 1 0 $X=142370 $Y=136000
X8536 3 1 470 384 DLY1JI3VX1 $T=143360 114240 1 0 $X=142930 $Y=109120
X8537 3 1 372 386 DLY1JI3VX1 $T=143920 51520 1 0 $X=143490 $Y=46400
X8538 3 1 1342 392 DLY1JI3VX1 $T=145040 176960 0 0 $X=144610 $Y=176320
X8539 3 1 398 850 DLY1JI3VX1 $T=145600 168000 1 0 $X=145170 $Y=162880
X8540 3 1 1228 399 DLY1JI3VX1 $T=150640 51520 1 0 $X=150210 $Y=46400
X8541 3 1 429 1171 DLY1JI3VX1 $T=150640 176960 0 0 $X=150210 $Y=176320
X8542 3 1 376 57 DLY1JI3VX1 $T=151200 168000 1 0 $X=150770 $Y=162880
X8543 3 1 1077 407 DLY1JI3VX1 $T=154000 123200 0 0 $X=153570 $Y=122560
X8544 3 1 444 408 DLY1JI3VX1 $T=154000 141120 1 0 $X=153570 $Y=136000
X8545 3 1 58 411 DLY1JI3VX1 $T=155120 150080 1 0 $X=154690 $Y=144960
X8546 3 1 402 1069 DLY1JI3VX1 $T=156240 51520 1 0 $X=155810 $Y=46400
X8547 3 1 865 1071 DLY1JI3VX1 $T=159040 168000 0 0 $X=158610 $Y=167360
X8548 3 1 412 421 DLY1JI3VX1 $T=160720 42560 1 0 $X=160290 $Y=37440
X8549 3 1 1232 862 DLY1JI3VX1 $T=164080 159040 1 0 $X=163650 $Y=153920
X8550 3 1 499 1305 DLY1JI3VX1 $T=164080 221760 1 0 $X=163650 $Y=216640
X8551 3 1 1346 864 DLY1JI3VX1 $T=166880 42560 1 0 $X=166450 $Y=37440
X8552 3 1 64 431 DLY1JI3VX1 $T=168000 78400 1 0 $X=167570 $Y=73280
X8553 3 1 423 432 DLY1JI3VX1 $T=168560 87360 1 0 $X=168130 $Y=82240
X8554 3 1 437 68 DLY1JI3VX1 $T=172480 42560 1 0 $X=172050 $Y=37440
X8555 3 1 469 85 DLY1JI3VX1 $T=183120 24640 1 180 $X=177090 $Y=24000
X8556 3 1 1235 450 DLY1JI3VX1 $T=178640 60480 1 0 $X=178210 $Y=55360
X8557 3 1 871 459 DLY1JI3VX1 $T=182560 150080 1 0 $X=182130 $Y=144960
X8558 3 1 1080 462 DLY1JI3VX1 $T=184240 194880 1 0 $X=183810 $Y=189760
X8559 3 1 1306 467 DLY1JI3VX1 $T=189280 33600 1 0 $X=188850 $Y=28480
X8560 3 1 466 468 DLY1JI3VX1 $T=189280 60480 1 0 $X=188850 $Y=55360
X8561 3 1 1307 1081 DLY1JI3VX1 $T=196000 78400 0 180 $X=189970 $Y=73280
X8562 3 1 964 875 DLY1JI3VX1 $T=194880 33600 1 0 $X=194450 $Y=28480
X8563 3 1 471 877 DLY1JI3VX1 $T=197680 141120 0 0 $X=197250 $Y=140480
X8564 3 1 81 476 DLY1JI3VX1 $T=199360 221760 1 0 $X=198930 $Y=216640
X8565 3 1 512 93 DLY1JI3VX1 $T=205520 60480 1 180 $X=199490 $Y=59840
X8566 3 1 881 82 DLY1JI3VX1 $T=203280 141120 0 0 $X=202850 $Y=140480
X8567 3 1 491 1310 DLY1JI3VX1 $T=211120 60480 1 180 $X=205090 $Y=59840
X8568 3 1 487 1363 DLY1JI3VX1 $T=211120 87360 0 180 $X=205090 $Y=82240
X8569 3 1 492 1176 DLY1JI3VX1 $T=211120 185920 0 180 $X=205090 $Y=180800
X8570 3 1 92 89 DLY1JI3VX1 $T=218960 176960 0 0 $X=218530 $Y=176320
X8571 3 1 513 91 DLY1JI3VX1 $T=225120 87360 0 180 $X=219090 $Y=82240
X8572 3 1 1242 505 DLY1JI3VX1 $T=230720 87360 0 180 $X=224690 $Y=82240
X8573 3 1 1243 90 DLY1JI3VX1 $T=235200 33600 0 180 $X=229170 $Y=28480
X8574 3 1 1096 519 DLY1JI3VX1 $T=230720 87360 1 0 $X=230290 $Y=82240
X8575 3 1 554 106 DLY1JI3VX1 $T=238000 87360 1 0 $X=237570 $Y=82240
X8576 3 1 114 544 DLY1JI3VX1 $T=240800 24640 0 0 $X=240370 $Y=24000
X8577 3 1 109 597 DLY1JI3VX1 $T=244160 168000 0 0 $X=243730 $Y=167360
X8578 3 1 540 550 DLY1JI3VX1 $T=244160 176960 1 0 $X=243730 $Y=171840
X8579 3 1 565 109 DLY1JI3VX1 $T=244720 159040 0 0 $X=244290 $Y=158400
X8580 3 1 548 557 DLY1JI3VX1 $T=248080 60480 0 0 $X=247650 $Y=59840
X8581 3 1 1248 563 DLY1JI3VX1 $T=250320 33600 1 0 $X=249890 $Y=28480
X8582 3 1 1178 115 DLY1JI3VX1 $T=251440 176960 1 0 $X=251010 $Y=171840
X8583 3 1 558 118 DLY1JI3VX1 $T=253680 60480 0 0 $X=253250 $Y=59840
X8584 3 1 1251 967 DLY1JI3VX1 $T=257040 176960 0 0 $X=256610 $Y=176320
X8585 3 1 1356 576 DLY1JI3VX1 $T=259840 42560 0 0 $X=259410 $Y=41920
X8586 3 1 610 594 DLY1JI3VX1 $T=262080 60480 0 0 $X=261650 $Y=59840
X8587 3 1 1252 120 DLY1JI3VX1 $T=265440 42560 0 0 $X=265010 $Y=41920
X8588 3 1 903 590 DLY1JI3VX1 $T=267680 176960 0 0 $X=267250 $Y=176320
X8589 3 1 588 905 DLY1JI3VX1 $T=271600 42560 0 0 $X=271170 $Y=41920
X8590 3 1 907 606 DLY1JI3VX1 $T=277200 42560 0 0 $X=276770 $Y=41920
X8591 3 1 909 613 DLY1JI3VX1 $T=282800 60480 0 0 $X=282370 $Y=59840
X8592 3 1 1257 911 DLY1JI3VX1 $T=283360 176960 0 0 $X=282930 $Y=176320
X8593 3 1 614 626 DLY1JI3VX1 $T=288400 60480 0 0 $X=287970 $Y=59840
X8594 3 1 616 628 DLY1JI3VX1 $T=288960 176960 0 0 $X=288530 $Y=176320
X8595 3 1 640 639 DLY1JI3VX1 $T=294560 60480 0 0 $X=294130 $Y=59840
X8596 3 1 1322 646 DLY1JI3VX1 $T=300160 42560 0 0 $X=299730 $Y=41920
X8597 3 1 1264 133 DLY1JI3VX1 $T=300160 60480 1 0 $X=299730 $Y=55360
X8598 3 1 113 648 DLY1JI3VX1 $T=302400 221760 1 0 $X=301970 $Y=216640
X8599 3 1 918 657 DLY1JI3VX1 $T=304080 87360 0 0 $X=303650 $Y=86720
X8600 3 1 655 1190 DLY1JI3VX1 $T=311360 60480 0 180 $X=305330 $Y=55360
X8601 3 1 647 664 DLY1JI3VX1 $T=306320 168000 0 0 $X=305890 $Y=167360
X8602 3 1 1268 671 DLY1JI3VX1 $T=309680 87360 1 0 $X=309250 $Y=82240
X8603 3 1 675 1359 DLY1JI3VX1 $T=316960 60480 0 180 $X=310930 $Y=55360
X8604 3 1 140 922 DLY1JI3VX1 $T=316960 150080 0 180 $X=310930 $Y=144960
X8605 3 1 141 1192 DLY1JI3VX1 $T=316960 150080 1 180 $X=310930 $Y=149440
X8606 3 1 692 145 DLY1JI3VX1 $T=324800 78400 0 0 $X=324370 $Y=77760
X8607 3 1 694 151 DLY1JI3VX1 $T=324800 105280 0 0 $X=324370 $Y=104640
X8608 3 1 1140 695 DLY1JI3VX1 $T=330400 51520 1 0 $X=329970 $Y=46400
X8609 3 1 1273 1148 DLY1JI3VX1 $T=334880 60480 1 0 $X=334450 $Y=55360
X8610 3 1 1380 705 DLY1JI3VX1 $T=334880 168000 1 0 $X=334450 $Y=162880
X8611 3 1 734 1194 DLY1JI3VX1 $T=340480 168000 1 0 $X=340050 $Y=162880
X8612 3 1 1327 1328 DLY1JI3VX1 $T=341040 60480 1 0 $X=340610 $Y=55360
X8613 3 1 1280 716 DLY1JI3VX1 $T=346640 60480 1 0 $X=346210 $Y=55360
X8614 3 1 1329 950 DLY1JI3VX1 $T=350000 150080 0 0 $X=349570 $Y=149440
X8615 3 1 1285 722 DLY1JI3VX1 $T=351680 42560 0 0 $X=351250 $Y=41920
X8616 3 1 731 723 DLY1JI3VX1 $T=351680 51520 1 0 $X=351250 $Y=46400
X8617 3 1 1286 725 DLY1JI3VX1 $T=352240 60480 1 0 $X=351810 $Y=55360
X8618 3 1 732 733 DLY1JI3VX1 $T=355600 150080 0 0 $X=355170 $Y=149440
X8619 3 1 954 738 DLY1JI3VX1 $T=358400 176960 0 0 $X=357970 $Y=176320
X8620 3 1 741 171 DLY1JI3VX1 $T=367360 60480 0 0 $X=366930 $Y=59840
X8621 3 1 1331 747 DLY1JI3VX1 $T=367920 51520 0 0 $X=367490 $Y=50880
X8622 3 1 955 748 DLY1JI3VX1 $T=373520 51520 0 0 $X=373090 $Y=50880
X8623 3 1 956 749 DLY1JI3VX1 $T=373520 60480 0 0 $X=373090 $Y=59840
X8624 3 1 1158 750 DLY1JI3VX1 $T=373520 176960 1 0 $X=373090 $Y=171840
X8625 3 1 174 751 DLY1JI3VX1 $T=374080 33600 1 0 $X=373650 $Y=28480
X8626 3 1 1291 757 DLY1JI3VX1 $T=379120 42560 1 0 $X=378690 $Y=37440
X8627 3 1 1293 758 DLY1JI3VX1 $T=379120 42560 0 0 $X=378690 $Y=41920
X8628 3 1 1292 759 DLY1JI3VX1 $T=379120 168000 1 0 $X=378690 $Y=162880
X8629 3 1 1397 404 1222 down_switches<21> ON21JI3VX4 $T=114800 24640 1 0 $X=114370 $Y=19520
X8630 3 1 1049 404 1225 down_switches<23> ON21JI3VX4 $T=124320 24640 1 0 $X=123890 $Y=19520
X8631 3 1 838 404 837 down_switches<20> ON21JI3VX4 $T=132720 24640 1 0 $X=132290 $Y=19520
X8632 3 1 849 404 1227 down_switches<22> ON21JI3VX4 $T=150080 24640 0 180 $X=141250 $Y=19520
X8633 3 1 845 404 962 down_switches<19> ON21JI3VX4 $T=146160 33600 1 0 $X=145730 $Y=28480
X8634 3 1 1062 404 1230 down_switches<18> ON21JI3VX4 $T=159040 24640 0 180 $X=150210 $Y=19520
X8635 3 1 1072 404 1233 down_switches<17> ON21JI3VX4 $T=168000 24640 0 180 $X=159170 $Y=19520
X8636 3 1 867 404 430 down_switches<16> ON21JI3VX4 $T=176400 24640 0 180 $X=167570 $Y=19520
X8637 3 1 1398 404 1076 down_switches<15> ON21JI3VX4 $T=182000 33600 0 180 $X=173170 $Y=28480
X8638 3 1 1399 404 1078 down_switches<14> ON21JI3VX4 $T=185360 24640 0 180 $X=176530 $Y=19520
X8639 3 1 1400 404 1369 down_switches<24> ON21JI3VX4 $T=194880 33600 1 180 $X=186050 $Y=32960
X8640 3 1 1401 404 1083 down_switches<13> ON21JI3VX4 $T=197680 24640 0 180 $X=188850 $Y=19520
X8641 3 1 884 404 1312 down_switches<26> ON21JI3VX4 $T=204400 24640 1 0 $X=203970 $Y=19520
X8642 3 1 1309 404 1087 down_switches<25> ON21JI3VX4 $T=204960 33600 1 0 $X=204530 $Y=28480
X8643 3 1 1090 404 1089 down_switches<27> ON21JI3VX4 $T=225120 33600 1 180 $X=216290 $Y=32960
X8644 3 1 1095 404 1240 down_switches<29> ON21JI3VX4 $T=228480 24640 0 180 $X=219650 $Y=19520
X8645 3 1 1402 404 1247 down_switches<30> ON21JI3VX4 $T=246960 33600 0 180 $X=238130 $Y=28480
X8646 3 1 899 404 1103 down_switches<28> ON21JI3VX4 $T=253120 33600 1 180 $X=244290 $Y=32960
X8647 3 1 1318 404 1253 down_switches<31> ON21JI3VX4 $T=270480 33600 0 180 $X=261650 $Y=28480
X8648 3 1 1255 404 1111 down_switches<12> ON21JI3VX4 $T=273840 24640 1 180 $X=265010 $Y=24000
X8649 3 1 1403 404 1320 down_switches<2> ON21JI3VX4 $T=283920 33600 0 180 $X=275090 $Y=28480
X8650 3 1 1260 404 1259 down_switches<3> ON21JI3VX4 $T=291200 33600 1 180 $X=282370 $Y=32960
X8651 3 1 914 404 1262 down_switches<0> ON21JI3VX4 $T=301840 33600 0 180 $X=293010 $Y=28480
X8652 3 1 921 404 1265 down_switches<11> ON21JI3VX4 $T=309120 24640 1 180 $X=300290 $Y=24000
X8653 3 1 1404 404 1378 down_switches<1> ON21JI3VX4 $T=310800 42560 1 0 $X=310370 $Y=37440
X8654 3 1 927 404 147 down_switches<10> ON21JI3VX4 $T=310800 42560 0 0 $X=310370 $Y=41920
X8655 3 1 1405 404 969 down_switches<4> ON21JI3VX4 $T=331520 33600 0 180 $X=322690 $Y=28480
X8656 3 1 1406 404 1379 down_switches<5> ON21JI3VX4 $T=337120 24640 0 180 $X=328290 $Y=19520
X8657 3 1 1147 404 1326 down_switches<9> ON21JI3VX4 $T=341040 33600 1 180 $X=332210 $Y=32960
X8658 3 1 949 404 1282 down_switches<8> ON21JI3VX4 $T=351680 33600 1 180 $X=342850 $Y=32960
X8659 3 1 1157 404 735 down_switches<6> ON21JI3VX4 $T=366240 24640 0 180 $X=357410 $Y=19520
X8660 3 1 1407 404 1289 down_switches<7> ON21JI3VX4 $T=367920 33600 0 180 $X=359090 $Y=28480
X8661 3 1 53 434 INJI3VX6 $T=176960 168000 1 0 $X=176530 $Y=162880
X8662 3 1 191 1408 186 979 NA3I1JI3VX1 $T=29680 60480 0 0 $X=29250 $Y=59840
X8663 3 1 13 1409 244 193 NA3I1JI3VX1 $T=56000 33600 1 180 $X=51650 $Y=32960
X8664 3 1 55 1362 785 244 NA3I1JI3VX1 $T=70000 33600 1 180 $X=65650 $Y=32960
X8665 3 1 821 812 814 813 NA3I1JI3VX1 $T=90160 194880 0 180 $X=85810 $Y=189760
X8666 3 1 100 1094 507 86 NA3I1JI3VX1 $T=227360 194880 0 0 $X=226930 $Y=194240
X8667 3 1 1094 1410 520 533 NA3I1JI3VX1 $T=236320 203840 1 0 $X=235890 $Y=198720
X8668 3 1 630 1395 624 627 NA3I1JI3VX1 $T=283360 212800 0 180 $X=279010 $Y=207680
X8669 3 1 668 pulse_active BUJI3VX8 $T=63840 24640 1 180 $X=55010 $Y=24000
X8670 3 1 1008 DAC<5> BUJI3VX8 $T=61600 24640 1 0 $X=61170 $Y=19520
X8671 3 1 1016 DAC<4> BUJI3VX8 $T=70560 24640 1 0 $X=70130 $Y=19520
X8672 3 1 1381 DAC<3> BUJI3VX8 $T=73360 24640 0 0 $X=72930 $Y=24000
X8673 3 1 1029 DAC<2> BUJI3VX8 $T=79520 24640 1 0 $X=79090 $Y=19520
X8674 3 1 1033 DAC<1> BUJI3VX8 $T=83440 24640 0 0 $X=83010 $Y=24000
X8675 3 1 1043 DAC<0> BUJI3VX8 $T=97440 24640 0 180 $X=88610 $Y=19520
X8676 3 1 66 4 BUJI3VX8 $T=173040 168000 1 180 $X=164210 $Y=167360
X8677 3 1 66 14 BUJI3VX8 $T=182560 78400 0 180 $X=173730 $Y=73280
X8678 3 1 66 111 BUJI3VX8 $T=190400 168000 0 180 $X=181570 $Y=162880
X8679 3 1 66 105 BUJI3VX8 $T=193760 87360 1 0 $X=193330 $Y=82240
X8680 3 1 180 763 4 182 DFRRQJI3VX1 $T=24080 123200 0 0 $X=23650 $Y=122560
X8681 3 1 180 176 4 179 DFRRQJI3VX1 $T=24080 141120 1 0 $X=23650 $Y=136000
X8682 3 1 180 177 4 5 DFRRQJI3VX1 $T=24080 141120 0 0 $X=23650 $Y=140480
X8683 3 1 180 1294 14 204 DFRRQJI3VX1 $T=24640 96320 0 0 $X=24210 $Y=95680
X8684 3 1 180 187 4 197 DFRRQJI3VX1 $T=24640 159040 1 0 $X=24210 $Y=153920
X8685 3 1 180 178 4 184 DFRRQJI3VX1 $T=24640 176960 1 0 $X=24210 $Y=171840
X8686 3 1 180 1332 14 13 DFRRQJI3VX1 $T=25200 33600 0 0 $X=24770 $Y=32960
X8687 3 1 180 190 14 10 DFRRQJI3VX1 $T=25200 42560 1 0 $X=24770 $Y=37440
X8688 3 1 180 1364 14 979 DFRRQJI3VX1 $T=25200 51520 0 0 $X=24770 $Y=50880
X8689 3 1 180 976 14 186 DFRRQJI3VX1 $T=25200 78400 1 0 $X=24770 $Y=73280
X8690 3 1 185 188 4 218 DFRRQJI3VX1 $T=25200 185920 1 0 $X=24770 $Y=180800
X8691 3 1 185 189 4 228 DFRRQJI3VX1 $T=25200 185920 0 0 $X=24770 $Y=185280
X8692 3 1 180 1202 14 984 DFRRQJI3VX1 $T=25760 87360 1 0 $X=25330 $Y=82240
X8693 3 1 180 181 14 8 DFRRQJI3VX1 $T=25760 96320 1 0 $X=25330 $Y=91200
X8694 3 1 185 762 4 9 DFRRQJI3VX1 $T=26320 194880 0 0 $X=25890 $Y=194240
X8695 3 1 185 977 4 227 DFRRQJI3VX1 $T=27440 212800 1 0 $X=27010 $Y=207680
X8696 3 1 180 988 4 11 DFRRQJI3VX1 $T=39200 132160 1 0 $X=38770 $Y=127040
X8697 3 1 180 989 4 20 DFRRQJI3VX1 $T=39760 132160 0 0 $X=39330 $Y=131520
X8698 3 1 180 769 4 198 DFRRQJI3VX1 $T=39760 141120 1 0 $X=39330 $Y=136000
X8699 3 1 185 776 4 201 DFRRQJI3VX1 $T=54880 168000 1 180 $X=39330 $Y=167360
X8700 3 1 180 214 14 196 DFRRQJI3VX1 $T=59360 87360 0 180 $X=43810 $Y=82240
X8701 3 1 185 1335 4 199 DFRRQJI3VX1 $T=44240 212800 1 0 $X=43810 $Y=207680
X8702 3 1 185 207 4 1007 DFRRQJI3VX1 $T=45360 212800 0 0 $X=44930 $Y=212160
X8703 3 1 180 1000 14 1010 DFRRQJI3VX1 $T=48160 78400 0 0 $X=47730 $Y=77760
X8704 3 1 180 220 14 222 DFRRQJI3VX1 $T=48720 69440 0 0 $X=48290 $Y=68800
X8705 3 1 180 19 14 1215 DFRRQJI3VX1 $T=48720 78400 1 0 $X=48290 $Y=73280
X8706 3 1 180 246 4 1209 DFRRQJI3VX1 $T=68320 159040 1 180 $X=52770 $Y=158400
X8707 3 1 180 787 4 237 DFRRQJI3VX1 $T=53760 159040 1 0 $X=53330 $Y=153920
X8708 3 1 180 223 4 794 DFRRQJI3VX1 $T=53760 168000 1 0 $X=53330 $Y=162880
X8709 3 1 180 1298 4 236 DFRRQJI3VX1 $T=54880 168000 0 0 $X=54450 $Y=167360
X8710 3 1 180 1214 4 782 DFRRQJI3VX1 $T=70560 132160 0 180 $X=55010 $Y=127040
X8711 3 1 180 243 4 795 DFRRQJI3VX1 $T=55440 141120 1 0 $X=55010 $Y=136000
X8712 3 1 180 238 4 256 DFRRQJI3VX1 $T=56560 114240 1 0 $X=56130 $Y=109120
X8713 3 1 180 226 4 793 DFRRQJI3VX1 $T=56560 123200 0 0 $X=56130 $Y=122560
X8714 3 1 180 797 14 55 DFRRQJI3VX1 $T=76160 51520 0 180 $X=60610 $Y=46400
X8715 3 1 180 258 14 217 DFRRQJI3VX1 $T=76720 51520 1 180 $X=61170 $Y=50880
X8716 3 1 180 245 14 16 DFRRQJI3VX1 $T=76720 60480 0 180 $X=61170 $Y=55360
X8717 3 1 185 1011 4 247 DFRRQJI3VX1 $T=61600 212800 0 0 $X=61170 $Y=212160
X8718 3 1 185 1018 4 232 DFRRQJI3VX1 $T=76720 221760 0 180 $X=61170 $Y=216640
X8719 3 1 180 251 14 248 DFRRQJI3VX1 $T=77280 60480 1 180 $X=61730 $Y=59840
X8720 3 1 180 287 14 241 DFRRQJI3VX1 $T=77840 69440 0 180 $X=62290 $Y=64320
X8721 3 1 180 1012 14 253 DFRRQJI3VX1 $T=63840 78400 0 0 $X=63410 $Y=77760
X8722 3 1 180 1014 14 257 DFRRQJI3VX1 $T=63840 87360 1 0 $X=63410 $Y=82240
X8723 3 1 180 288 14 224 DFRRQJI3VX1 $T=79520 69440 1 180 $X=63970 $Y=68800
X8724 3 1 180 255 4 263 DFRRQJI3VX1 $T=69440 150080 0 0 $X=69010 $Y=149440
X8725 3 1 180 30 4 230 DFRRQJI3VX1 $T=84560 159040 0 180 $X=69010 $Y=153920
X8726 3 1 180 804 4 234 DFRRQJI3VX1 $T=84560 168000 0 180 $X=69010 $Y=162880
X8727 3 1 180 271 4 278 DFRRQJI3VX1 $T=84560 176960 0 180 $X=69010 $Y=171840
X8728 3 1 180 264 4 1015 DFRRQJI3VX1 $T=85120 168000 1 180 $X=69570 $Y=167360
X8729 3 1 180 267 14 316 DFRRQJI3VX1 $T=77840 42560 1 0 $X=77410 $Y=37440
X8730 3 1 180 289 14 301 DFRRQJI3VX1 $T=77840 42560 0 0 $X=77410 $Y=41920
X8731 3 1 180 28 14 262 DFRRQJI3VX1 $T=92960 51520 0 180 $X=77410 $Y=46400
X8732 3 1 185 268 4 265 DFRRQJI3VX1 $T=93520 212800 1 180 $X=77970 $Y=212160
X8733 3 1 185 1032 4 282 DFRRQJI3VX1 $T=78400 221760 1 0 $X=77970 $Y=216640
X8734 3 1 180 1036 14 822 DFRRQJI3VX1 $T=79520 87360 1 0 $X=79090 $Y=82240
X8735 3 1 180 285 4 31 DFRRQJI3VX1 $T=99680 150080 0 180 $X=84130 $Y=144960
X8736 3 1 180 297 4 810 DFRRQJI3VX1 $T=100240 150080 1 180 $X=84690 $Y=149440
X8737 3 1 180 298 4 1034 DFRRQJI3VX1 $T=100240 159040 0 180 $X=84690 $Y=153920
X8738 3 1 180 299 4 293 DFRRQJI3VX1 $T=85680 159040 0 0 $X=85250 $Y=158400
X8739 3 1 180 304 4 811 DFRRQJI3VX1 $T=100800 168000 0 180 $X=85250 $Y=162880
X8740 3 1 180 1367 4 274 DFRRQJI3VX1 $T=100800 176960 0 180 $X=85250 $Y=171840
X8741 3 1 180 39 4 242 DFRRQJI3VX1 $T=101360 168000 1 180 $X=85810 $Y=167360
X8742 3 1 180 290 14 270 DFRRQJI3VX1 $T=104720 114240 1 180 $X=89170 $Y=113600
X8743 3 1 180 291 14 26 DFRRQJI3VX1 $T=104720 123200 0 180 $X=89170 $Y=118080
X8744 3 1 53 1338 14 826 DFRRQJI3VX1 $T=109200 33600 0 180 $X=93650 $Y=28480
X8745 3 1 53 300 14 1166 DFRRQJI3VX1 $T=109200 33600 1 180 $X=93650 $Y=32960
X8746 3 1 53 1039 14 37 DFRRQJI3VX1 $T=109760 42560 0 180 $X=94210 $Y=37440
X8747 3 1 180 295 14 1044 DFRRQJI3VX1 $T=109760 51520 0 180 $X=94210 $Y=46400
X8748 3 1 180 42 14 215 DFRRQJI3VX1 $T=109760 78400 1 180 $X=94210 $Y=77760
X8749 3 1 180 302 14 225 DFRRQJI3VX1 $T=109760 87360 1 180 $X=94210 $Y=86720
X8750 3 1 180 309 14 280 DFRRQJI3VX1 $T=109760 96320 0 180 $X=94210 $Y=91200
X8751 3 1 180 310 14 33 DFRRQJI3VX1 $T=110320 96320 1 180 $X=94770 $Y=95680
X8752 3 1 180 827 14 818 DFRRQJI3VX1 $T=110320 114240 0 180 $X=94770 $Y=109120
X8753 3 1 185 1340 4 38 DFRRQJI3VX1 $T=110320 203840 0 180 $X=94770 $Y=198720
X8754 3 1 185 1339 4 308 DFRRQJI3VX1 $T=110320 212800 0 180 $X=94770 $Y=207680
X8755 3 1 185 830 4 1041 DFRRQJI3VX1 $T=110320 221760 0 180 $X=94770 $Y=216640
X8756 3 1 53 344 4 321 DFRRQJI3VX1 $T=108080 168000 1 0 $X=107650 $Y=162880
X8757 3 1 53 47 4 1048 DFRRQJI3VX1 $T=108080 168000 0 0 $X=107650 $Y=167360
X8758 3 1 53 339 4 318 DFRRQJI3VX1 $T=108080 176960 0 0 $X=107650 $Y=176320
X8759 3 1 185 1223 4 319 DFRRQJI3VX1 $T=108080 203840 0 0 $X=107650 $Y=203200
X8760 3 1 185 320 4 833 DFRRQJI3VX1 $T=108080 212800 0 0 $X=107650 $Y=212160
X8761 3 1 53 832 14 323 DFRRQJI3VX1 $T=109760 105280 1 0 $X=109330 $Y=100160
X8762 3 1 53 364 14 325 DFRRQJI3VX1 $T=110880 96320 1 0 $X=110450 $Y=91200
X8763 3 1 53 334 14 326 DFRRQJI3VX1 $T=110880 105280 0 0 $X=110450 $Y=104640
X8764 3 1 53 305 14 835 DFRRQJI3VX1 $T=111440 33600 1 0 $X=111010 $Y=28480
X8765 3 1 53 315 14 374 DFRRQJI3VX1 $T=111440 33600 0 0 $X=111010 $Y=32960
X8766 3 1 53 306 14 327 DFRRQJI3VX1 $T=111440 42560 1 0 $X=111010 $Y=37440
X8767 3 1 53 340 14 328 DFRRQJI3VX1 $T=111440 42560 0 0 $X=111010 $Y=41920
X8768 3 1 53 341 14 347 DFRRQJI3VX1 $T=111440 51520 0 0 $X=111010 $Y=50880
X8769 3 1 53 380 14 329 DFRRQJI3VX1 $T=111440 87360 0 0 $X=111010 $Y=86720
X8770 3 1 53 342 14 324 DFRRQJI3VX1 $T=112000 51520 1 0 $X=111570 $Y=46400
X8771 3 1 53 317 14 986 DFRRQJI3VX1 $T=112560 114240 1 0 $X=112130 $Y=109120
X8772 3 1 53 335 4 834 DFRRQJI3VX1 $T=117600 185920 1 0 $X=117170 $Y=180800
X8773 3 1 53 349 4 51 DFRRQJI3VX1 $T=133280 176960 0 180 $X=117730 $Y=171840
X8774 3 1 185 360 4 369 DFRRQJI3VX1 $T=122640 221760 1 0 $X=122210 $Y=216640
X8775 3 1 53 391 4 376 DFRRQJI3VX1 $T=127120 168000 1 0 $X=126690 $Y=162880
X8776 3 1 53 337 4 1342 DFRRQJI3VX1 $T=127120 168000 0 0 $X=126690 $Y=167360
X8777 3 1 53 378 14 330 DFRRQJI3VX1 $T=143360 87360 1 180 $X=127810 $Y=86720
X8778 3 1 56 370 14 831 DFRRQJI3VX1 $T=143360 105280 0 180 $X=127810 $Y=100160
X8779 3 1 53 365 14 331 DFRRQJI3VX1 $T=143360 105280 1 180 $X=127810 $Y=104640
X8780 3 1 53 384 14 333 DFRRQJI3VX1 $T=143360 114240 0 180 $X=127810 $Y=109120
X8781 3 1 53 1069 14 354 DFRRQJI3VX1 $T=143920 42560 0 180 $X=128370 $Y=37440
X8782 3 1 53 356 14 389 DFRRQJI3VX1 $T=128800 42560 0 0 $X=128370 $Y=41920
X8783 3 1 53 386 14 385 DFRRQJI3VX1 $T=128800 51520 1 0 $X=128370 $Y=46400
X8784 3 1 53 357 14 1056 DFRRQJI3VX1 $T=128800 51520 0 0 $X=128370 $Y=50880
X8785 3 1 53 367 4 1037 DFRRQJI3VX1 $T=143920 123200 0 180 $X=128370 $Y=118080
X8786 3 1 53 392 4 350 DFRRQJI3VX1 $T=145040 176960 1 180 $X=129490 $Y=176320
X8787 3 1 53 358 14 402 DFRRQJI3VX1 $T=133280 60480 1 0 $X=132850 $Y=55360
X8788 3 1 53 375 14 372 DFRRQJI3VX1 $T=148400 60480 1 180 $X=132850 $Y=59840
X8789 3 1 56 352 14 381 DFRRQJI3VX1 $T=133280 69440 1 0 $X=132850 $Y=64320
X8790 3 1 53 382 4 345 DFRRQJI3VX1 $T=148400 159040 0 180 $X=132850 $Y=153920
X8791 3 1 185 1343 4 395 DFRRQJI3VX1 $T=138880 212800 0 0 $X=138450 $Y=212160
X8792 3 1 185 844 4 852 DFRRQJI3VX1 $T=138880 221760 1 0 $X=138450 $Y=216640
X8793 3 1 56 390 4 398 DFRRQJI3VX1 $T=139440 159040 0 0 $X=139010 $Y=158400
X8794 3 1 53 850 4 840 DFRRQJI3VX1 $T=155680 176960 0 180 $X=140130 $Y=171840
X8795 3 1 53 57 4 1055 DFRRQJI3VX1 $T=157360 168000 1 180 $X=141810 $Y=167360
X8796 3 1 56 406 4 366 DFRRQJI3VX1 $T=158480 105280 1 180 $X=142930 $Y=104640
X8797 3 1 56 1060 4 371 DFRRQJI3VX1 $T=159040 114240 1 180 $X=143490 $Y=113600
X8798 3 1 56 407 4 842 DFRRQJI3VX1 $T=159040 123200 0 180 $X=143490 $Y=118080
X8799 3 1 56 408 4 373 DFRRQJI3VX1 $T=159600 132160 1 180 $X=144050 $Y=131520
X8800 3 1 56 421 14 410 DFRRQJI3VX1 $T=145600 42560 1 0 $X=145170 $Y=37440
X8801 3 1 56 399 14 857 DFRRQJI3VX1 $T=145600 42560 0 0 $X=145170 $Y=41920
X8802 3 1 56 414 14 1346 DFRRQJI3VX1 $T=145600 51520 0 0 $X=145170 $Y=50880
X8803 3 1 56 411 4 379 DFRRQJI3VX1 $T=160720 150080 1 180 $X=145170 $Y=149440
X8804 3 1 56 418 14 1228 DFRRQJI3VX1 $T=163520 60480 0 180 $X=147970 $Y=55360
X8805 3 1 56 415 14 412 DFRRQJI3VX1 $T=163520 60480 1 180 $X=147970 $Y=59840
X8806 3 1 56 396 14 423 DFRRQJI3VX1 $T=148400 69440 1 0 $X=147970 $Y=64320
X8807 3 1 56 401 4 1232 DFRRQJI3VX1 $T=148400 159040 1 0 $X=147970 $Y=153920
X8808 3 1 185 1347 4 856 DFRRQJI3VX1 $T=170240 212800 1 180 $X=154690 $Y=212160
X8809 3 1 56 862 4 854 DFRRQJI3VX1 $T=170800 159040 1 180 $X=155250 $Y=158400
X8810 3 1 185 1066 4 426 DFRRQJI3VX1 $T=155680 212800 1 0 $X=155250 $Y=207680
X8811 3 1 53 1071 4 1063 DFRRQJI3VX1 $T=171360 176960 0 180 $X=155810 $Y=171840
X8812 3 1 53 1171 4 419 DFRRQJI3VX1 $T=171360 176960 1 180 $X=155810 $Y=176320
X8813 3 1 56 438 4 865 DFRRQJI3VX1 $T=156800 168000 1 0 $X=156370 $Y=162880
X8814 3 1 56 432 14 1068 DFRRQJI3VX1 $T=174160 33600 1 180 $X=158610 $Y=32960
X8815 3 1 56 864 14 425 DFRRQJI3VX1 $T=177520 42560 1 180 $X=161970 $Y=41920
X8816 3 1 71 431 14 869 DFRRQJI3VX1 $T=162960 51520 1 0 $X=162530 $Y=46400
X8817 3 1 56 68 14 61 DFRRQJI3VX1 $T=178080 51520 1 180 $X=162530 $Y=50880
X8818 3 1 56 450 14 1070 DFRRQJI3VX1 $T=178640 60480 0 180 $X=163090 $Y=55360
X8819 3 1 71 455 14 1235 DFRRQJI3VX1 $T=163520 60480 0 0 $X=163090 $Y=59840
X8820 3 1 71 454 14 437 DFRRQJI3VX1 $T=163520 69440 1 0 $X=163090 $Y=64320
X8821 3 1 56 456 14 64 DFRRQJI3VX1 $T=178640 69440 1 180 $X=163090 $Y=68800
X8822 3 1 185 445 111 442 DFRRQJI3VX1 $T=187040 212800 0 180 $X=171490 $Y=207680
X8823 3 1 185 1348 111 75 DFRRQJI3VX1 $T=171920 212800 0 0 $X=171490 $Y=212160
X8824 3 1 185 436 111 1079 DFRRQJI3VX1 $T=172480 203840 0 0 $X=172050 $Y=203200
X8825 3 1 56 74 111 427 DFRRQJI3VX1 $T=188160 159040 1 180 $X=172610 $Y=158400
X8826 3 1 56 449 111 429 DFRRQJI3VX1 $T=188160 168000 1 180 $X=172610 $Y=167360
X8827 3 1 56 459 111 1074 DFRRQJI3VX1 $T=188160 176960 0 180 $X=172610 $Y=171840
X8828 3 1 71 441 111 1080 DFRRQJI3VX1 $T=173040 176960 0 0 $X=172610 $Y=176320
X8829 3 1 185 462 111 439 DFRRQJI3VX1 $T=188160 185920 0 180 $X=172610 $Y=180800
X8830 3 1 71 875 14 870 DFRRQJI3VX1 $T=194320 42560 1 180 $X=178770 $Y=41920
X8831 3 1 71 67 14 964 DFRRQJI3VX1 $T=179200 69440 1 0 $X=178770 $Y=64320
X8832 3 1 71 467 14 457 DFRRQJI3VX1 $T=194880 51520 0 180 $X=179330 $Y=46400
X8833 3 1 71 468 14 453 DFRRQJI3VX1 $T=194880 51520 1 180 $X=179330 $Y=50880
X8834 3 1 71 1174 14 466 DFRRQJI3VX1 $T=179760 60480 0 0 $X=179330 $Y=59840
X8835 3 1 71 463 14 1306 DFRRQJI3VX1 $T=179760 69440 0 0 $X=179330 $Y=68800
X8836 3 1 71 591 14 440 DFRRQJI3VX1 $T=197680 114240 0 180 $X=182130 $Y=109120
X8837 3 1 71 521 14 443 DFRRQJI3VX1 $T=197680 114240 1 180 $X=182130 $Y=113600
X8838 3 1 71 564 14 1077 DFRRQJI3VX1 $T=197680 123200 1 180 $X=182130 $Y=122560
X8839 3 1 71 538 111 444 DFRRQJI3VX1 $T=197680 132160 1 180 $X=182130 $Y=131520
X8840 3 1 71 502 111 58 DFRRQJI3VX1 $T=197680 141120 1 180 $X=182130 $Y=140480
X8841 3 1 185 475 111 474 DFRRQJI3VX1 $T=188160 212800 1 0 $X=187730 $Y=207680
X8842 3 1 185 1370 111 473 DFRRQJI3VX1 $T=188720 203840 0 0 $X=188290 $Y=203200
X8843 3 1 71 476 111 461 DFRRQJI3VX1 $T=204960 185920 0 180 $X=189410 $Y=180800
X8844 3 1 71 481 111 881 DFRRQJI3VX1 $T=190960 150080 1 0 $X=190530 $Y=144960
X8845 3 1 71 529 111 871 DFRRQJI3VX1 $T=206080 168000 0 180 $X=190530 $Y=162880
X8846 3 1 71 530 111 81 DFRRQJI3VX1 $T=206080 168000 1 180 $X=190530 $Y=167360
X8847 3 1 71 82 111 872 DFRRQJI3VX1 $T=206080 176960 0 180 $X=190530 $Y=171840
X8848 3 1 71 501 111 446 DFRRQJI3VX1 $T=206640 141120 0 180 $X=191090 $Y=136000
X8849 3 1 71 458 111 471 DFRRQJI3VX1 $T=206640 159040 1 180 $X=191090 $Y=158400
X8850 3 1 71 877 111 965 DFRRQJI3VX1 $T=191520 176960 0 0 $X=191090 $Y=176320
X8851 3 1 71 479 14 469 DFRRQJI3VX1 $T=211120 69440 0 180 $X=195570 $Y=64320
X8852 3 1 71 87 14 1307 DFRRQJI3VX1 $T=211120 78400 0 180 $X=195570 $Y=73280
X8853 3 1 71 85 14 1308 DFRRQJI3VX1 $T=211680 42560 1 180 $X=196130 $Y=41920
X8854 3 1 71 1310 14 880 DFRRQJI3VX1 $T=211680 51520 0 180 $X=196130 $Y=46400
X8855 3 1 71 1175 14 491 DFRRQJI3VX1 $T=211680 51520 1 180 $X=196130 $Y=50880
X8856 3 1 71 1081 14 874 DFRRQJI3VX1 $T=211680 60480 0 180 $X=196130 $Y=55360
X8857 3 1 71 1363 14 873 DFRRQJI3VX1 $T=211680 69440 1 180 $X=196130 $Y=68800
X8858 3 1 71 84 14 487 DFRRQJI3VX1 $T=211680 78400 1 180 $X=196130 $Y=77760
X8859 3 1 71 531 14 465 DFRRQJI3VX1 $T=212240 105280 0 180 $X=196690 $Y=100160
X8860 3 1 71 532 14 470 DFRRQJI3VX1 $T=213920 114240 0 180 $X=198370 $Y=109120
X8861 3 1 71 527 14 472 DFRRQJI3VX1 $T=213920 114240 1 180 $X=198370 $Y=113600
X8862 3 1 185 883 111 1084 DFRRQJI3VX1 $T=215040 212800 1 180 $X=199490 $Y=212160
X8863 3 1 518 505 105 101 DFRRQJI3VX1 $T=213920 51520 0 0 $X=213490 $Y=50880
X8864 3 1 518 88 111 92 DFRRQJI3VX1 $T=213920 168000 1 0 $X=213490 $Y=162880
X8865 3 1 71 89 111 509 DFRRQJI3VX1 $T=213920 168000 0 0 $X=213490 $Y=167360
X8866 3 1 518 1176 111 98 DFRRQJI3VX1 $T=213920 176960 1 0 $X=213490 $Y=171840
X8867 3 1 108 524 111 492 DFRRQJI3VX1 $T=213920 185920 1 0 $X=213490 $Y=180800
X8868 3 1 108 1349 111 885 DFRRQJI3VX1 $T=213920 212800 1 0 $X=213490 $Y=207680
X8869 3 1 518 519 105 510 DFRRQJI3VX1 $T=214480 42560 0 0 $X=214050 $Y=41920
X8870 3 1 518 90 105 1092 DFRRQJI3VX1 $T=214480 51520 1 0 $X=214050 $Y=46400
X8871 3 1 518 91 105 511 DFRRQJI3VX1 $T=214480 60480 1 0 $X=214050 $Y=55360
X8872 3 1 518 93 105 887 DFRRQJI3VX1 $T=214480 60480 0 0 $X=214050 $Y=59840
X8873 3 1 518 96 105 1243 DFRRQJI3VX1 $T=214480 69440 1 0 $X=214050 $Y=64320
X8874 3 1 518 526 105 512 DFRRQJI3VX1 $T=214480 69440 0 0 $X=214050 $Y=68800
X8875 3 1 518 525 105 513 DFRRQJI3VX1 $T=214480 78400 1 0 $X=214050 $Y=73280
X8876 3 1 518 95 105 1242 DFRRQJI3VX1 $T=214480 78400 0 0 $X=214050 $Y=77760
X8877 3 1 108 886 111 507 DFRRQJI3VX1 $T=217840 212800 0 0 $X=217410 $Y=212160
X8878 3 1 108 552 111 1178 DFRRQJI3VX1 $T=226800 176960 0 0 $X=226370 $Y=176320
X8879 3 1 108 893 111 540 DFRRQJI3VX1 $T=244160 168000 1 180 $X=228610 $Y=167360
X8880 3 1 108 550 111 1101 DFRRQJI3VX1 $T=229040 176960 1 0 $X=228610 $Y=171840
X8881 3 1 108 537 111 520 DFRRQJI3VX1 $T=246400 212800 0 180 $X=230850 $Y=207680
X8882 3 1 518 569 105 1248 DFRRQJI3VX1 $T=231840 78400 1 0 $X=231410 $Y=73280
X8883 3 1 518 586 105 558 DFRRQJI3VX1 $T=231840 78400 0 0 $X=231410 $Y=77760
X8884 3 1 518 544 105 1098 DFRRQJI3VX1 $T=247520 42560 1 180 $X=231970 $Y=41920
X8885 3 1 518 563 105 889 DFRRQJI3VX1 $T=247520 51520 0 180 $X=231970 $Y=46400
X8886 3 1 518 557 105 543 DFRRQJI3VX1 $T=232400 51520 0 0 $X=231970 $Y=50880
X8887 3 1 518 118 105 1097 DFRRQJI3VX1 $T=247520 60480 0 180 $X=231970 $Y=55360
X8888 3 1 518 106 105 896 DFRRQJI3VX1 $T=232960 60480 0 0 $X=232530 $Y=59840
X8889 3 1 518 568 105 1096 DFRRQJI3VX1 $T=248080 69440 0 180 $X=232530 $Y=64320
X8890 3 1 518 102 105 548 DFRRQJI3VX1 $T=248080 69440 1 180 $X=232530 $Y=68800
X8891 3 1 108 546 111 522 DFRRQJI3VX1 $T=253680 194880 1 180 $X=238130 $Y=194240
X8892 3 1 108 562 111 542 DFRRQJI3VX1 $T=253680 203840 1 180 $X=238130 $Y=203200
X8893 3 1 108 967 111 99 DFRRQJI3VX1 $T=255920 185920 0 180 $X=240370 $Y=180800
X8894 3 1 108 110 111 1251 DFRRQJI3VX1 $T=241360 185920 0 0 $X=240930 $Y=185280
X8895 3 1 108 115 111 894 DFRRQJI3VX1 $T=257040 176960 1 180 $X=241490 $Y=176320
X8896 3 1 518 120 105 897 DFRRQJI3VX1 $T=265440 51520 0 180 $X=249890 $Y=46400
X8897 3 1 518 576 105 898 DFRRQJI3VX1 $T=265440 51520 1 180 $X=249890 $Y=50880
X8898 3 1 518 585 105 114 DFRRQJI3VX1 $T=265440 60480 0 180 $X=249890 $Y=55360
X8899 3 1 518 584 105 1356 DFRRQJI3VX1 $T=250320 69440 1 0 $X=249890 $Y=64320
X8900 3 1 518 587 105 1252 DFRRQJI3VX1 $T=250320 69440 0 0 $X=249890 $Y=68800
X8901 3 1 518 572 105 554 DFRRQJI3VX1 $T=267120 105280 0 180 $X=251570 $Y=100160
X8902 3 1 108 590 111 553 DFRRQJI3VX1 $T=273280 185920 1 180 $X=257730 $Y=185280
X8903 3 1 604 573 111 903 DFRRQJI3VX1 $T=258720 185920 1 0 $X=258290 $Y=180800
X8904 3 1 618 1112 116 1118 DFRRQJI3VX1 $T=266000 203840 0 0 $X=265570 $Y=203200
X8905 3 1 618 1254 116 603 DFRRQJI3VX1 $T=266000 212800 0 0 $X=265570 $Y=212160
X8906 3 1 108 123 105 909 DFRRQJI3VX1 $T=267120 105280 1 0 $X=266690 $Y=100160
X8907 3 1 518 905 105 595 DFRRQJI3VX1 $T=282800 51520 0 180 $X=267250 $Y=46400
X8908 3 1 518 606 105 902 DFRRQJI3VX1 $T=282800 51520 1 180 $X=267250 $Y=50880
X8909 3 1 518 615 105 907 DFRRQJI3VX1 $T=267680 60480 1 0 $X=267250 $Y=55360
X8910 3 1 518 626 105 582 DFRRQJI3VX1 $T=282800 60480 1 180 $X=267250 $Y=59840
X8911 3 1 518 613 105 124 DFRRQJI3VX1 $T=282800 69440 0 180 $X=267250 $Y=64320
X8912 3 1 518 619 105 588 DFRRQJI3VX1 $T=282800 69440 1 180 $X=267250 $Y=68800
X8913 3 1 518 594 105 1258 DFRRQJI3VX1 $T=269360 42560 1 0 $X=268930 $Y=37440
X8914 3 1 154 621 105 610 DFRRQJI3VX1 $T=272160 78400 1 0 $X=271730 $Y=73280
X8915 3 1 154 666 105 614 DFRRQJI3VX1 $T=292320 114240 1 180 $X=276770 $Y=113600
X8916 3 1 618 1119 116 624 DFRRQJI3VX1 $T=277200 194880 0 0 $X=276770 $Y=194240
X8917 3 1 633 911 111 1127 DFRRQJI3VX1 $T=279440 185920 1 0 $X=279010 $Y=180800
X8918 3 1 908 636 111 1257 DFRRQJI3VX1 $T=295120 176960 0 180 $X=279570 $Y=171840
X8919 3 1 618 634 116 630 DFRRQJI3VX1 $T=297920 203840 1 180 $X=282370 $Y=203200
X8920 3 1 1261 628 111 1128 DFRRQJI3VX1 $T=283920 168000 0 0 $X=283490 $Y=167360
X8921 3 1 618 1357 116 617 DFRRQJI3VX1 $T=299040 212800 1 180 $X=283490 $Y=212160
X8922 3 1 611 638 111 616 DFRRQJI3VX1 $T=299600 168000 0 180 $X=284050 $Y=162880
X8923 3 1 633 1122 111 912 DFRRQJI3VX1 $T=284480 185920 0 0 $X=284050 $Y=185280
X8924 3 1 518 646 105 1121 DFRRQJI3VX1 $T=300160 42560 1 180 $X=284610 $Y=41920
X8925 3 1 518 133 105 629 DFRRQJI3VX1 $T=300160 51520 0 180 $X=284610 $Y=46400
X8926 3 1 518 639 105 910 DFRRQJI3VX1 $T=300160 51520 1 180 $X=284610 $Y=50880
X8927 3 1 154 651 105 1322 DFRRQJI3VX1 $T=285040 60480 1 0 $X=284610 $Y=55360
X8928 3 1 154 656 105 1264 DFRRQJI3VX1 $T=285040 69440 1 0 $X=284610 $Y=64320
X8929 3 1 154 622 105 640 DFRRQJI3VX1 $T=285040 69440 0 0 $X=284610 $Y=68800
X8930 3 1 154 652 105 918 DFRRQJI3VX1 $T=294000 96320 0 0 $X=293570 $Y=95680
X8931 3 1 154 653 105 1268 DFRRQJI3VX1 $T=294000 105280 1 0 $X=293570 $Y=100160
X8932 3 1 154 671 105 637 DFRRQJI3VX1 $T=309680 87360 0 180 $X=294130 $Y=82240
X8933 3 1 154 657 105 1124 DFRRQJI3VX1 $T=309680 96320 0 180 $X=294130 $Y=91200
X8934 3 1 677 1129 111 1411 DFRRQJI3VX1 $T=297920 203840 1 0 $X=297490 $Y=198720
X8935 3 1 913 1358 111 662 DFRRQJI3VX1 $T=313600 203840 1 180 $X=298050 $Y=203200
X8936 3 1 919 136 111 647 DFRRQJI3VX1 $T=315840 159040 1 180 $X=300290 $Y=158400
X8937 3 1 1132 664 111 1133 DFRRQJI3VX1 $T=300720 168000 1 0 $X=300290 $Y=162880
X8938 3 1 154 1359 105 1130 DFRRQJI3VX1 $T=316960 51520 0 180 $X=301410 $Y=46400
X8939 3 1 154 1190 105 915 DFRRQJI3VX1 $T=316960 51520 1 180 $X=301410 $Y=50880
X8940 3 1 154 710 105 675 DFRRQJI3VX1 $T=316960 60480 1 180 $X=301410 $Y=59840
X8941 3 1 154 709 105 655 DFRRQJI3VX1 $T=316960 69440 0 180 $X=301410 $Y=64320
X8942 3 1 154 922 111 916 DFRRQJI3VX1 $T=317520 159040 0 180 $X=301970 $Y=153920
X8943 3 1 659 679 111 142 DFRRQJI3VX1 $T=322000 212800 0 180 $X=306450 $Y=207680
X8944 3 1 1267 144 111 665 DFRRQJI3VX1 $T=322000 212800 1 180 $X=306450 $Y=212160
X8945 3 1 154 695 105 157 DFRRQJI3VX1 $T=319760 51520 0 0 $X=319330 $Y=50880
X8946 3 1 154 1148 105 691 DFRRQJI3VX1 $T=319760 60480 1 0 $X=319330 $Y=55360
X8947 3 1 154 148 105 1273 DFRRQJI3VX1 $T=319760 60480 0 0 $X=319330 $Y=59840
X8948 3 1 154 711 105 1140 DFRRQJI3VX1 $T=319760 69440 1 0 $X=319330 $Y=64320
X8949 3 1 154 145 105 693 DFRRQJI3VX1 $T=319760 96320 1 0 $X=319330 $Y=91200
X8950 3 1 154 151 105 1135 DFRRQJI3VX1 $T=319760 96320 0 0 $X=319330 $Y=95680
X8951 3 1 154 683 105 692 DFRRQJI3VX1 $T=319760 105280 1 0 $X=319330 $Y=100160
X8952 3 1 154 681 105 694 DFRRQJI3VX1 $T=319760 114240 1 0 $X=319330 $Y=109120
X8953 3 1 154 712 111 140 DFRRQJI3VX1 $T=319760 141120 1 0 $X=319330 $Y=136000
X8954 3 1 154 149 111 141 DFRRQJI3VX1 $T=319760 141120 0 0 $X=319330 $Y=140480
X8955 3 1 154 1192 111 152 DFRRQJI3VX1 $T=319760 150080 0 0 $X=319330 $Y=149440
X8956 3 1 161 685 111 1380 DFRRQJI3VX1 $T=319760 159040 0 0 $X=319330 $Y=158400
X8957 3 1 700 705 111 931 DFRRQJI3VX1 $T=319760 168000 1 0 $X=319330 $Y=162880
X8958 3 1 161 721 111 1329 DFRRQJI3VX1 $T=334880 141120 0 0 $X=334450 $Y=140480
X8959 3 1 161 950 111 1274 DFRRQJI3VX1 $T=350000 150080 1 180 $X=334450 $Y=149440
X8960 3 1 154 722 105 1145 DFRRQJI3VX1 $T=351680 42560 1 180 $X=336130 $Y=41920
X8961 3 1 154 723 105 932 DFRRQJI3VX1 $T=351680 51520 0 180 $X=336130 $Y=46400
X8962 3 1 154 1328 105 1277 DFRRQJI3VX1 $T=351680 51520 1 180 $X=336130 $Y=50880
X8963 3 1 154 725 105 158 DFRRQJI3VX1 $T=351680 60480 1 180 $X=336130 $Y=59840
X8964 3 1 154 720 105 1286 DFRRQJI3VX1 $T=336560 105280 1 0 $X=336130 $Y=100160
X8965 3 1 154 716 105 938 DFRRQJI3VX1 $T=352240 69440 0 180 $X=336690 $Y=64320
X8966 3 1 154 708 105 1285 DFRRQJI3VX1 $T=337120 96320 0 0 $X=336690 $Y=95680
X8967 3 1 154 728 105 1327 DFRRQJI3VX1 $T=360080 69440 1 180 $X=344530 $Y=68800
X8968 3 1 154 724 105 1280 DFRRQJI3VX1 $T=360080 78400 0 180 $X=344530 $Y=73280
X8969 3 1 154 1156 105 731 DFRRQJI3VX1 $T=344960 87360 0 0 $X=344530 $Y=86720
X8970 3 1 161 733 111 713 DFRRQJI3VX1 $T=361200 159040 1 180 $X=345650 $Y=158400
X8971 3 1 161 1194 111 714 DFRRQJI3VX1 $T=361200 168000 0 180 $X=345650 $Y=162880
X8972 3 1 161 717 111 954 DFRRQJI3VX1 $T=346640 150080 1 0 $X=346210 $Y=144960
X8973 3 1 161 168 111 732 DFRRQJI3VX1 $T=346640 159040 1 0 $X=346210 $Y=153920
X8974 3 1 161 738 111 944 DFRRQJI3VX1 $T=361760 168000 1 180 $X=346210 $Y=167360
X8975 3 1 154 171 105 952 DFRRQJI3VX1 $T=367360 60480 1 180 $X=351810 $Y=59840
X8976 3 1 154 726 105 1331 DFRRQJI3VX1 $T=352240 69440 1 0 $X=351810 $Y=64320
X8977 3 1 1287 1200 111 727 DFRRQJI3VX1 $T=367360 203840 0 180 $X=351810 $Y=198720
X8978 3 1 154 747 105 160 DFRRQJI3VX1 $T=367920 51520 1 180 $X=352370 $Y=50880
X8979 3 1 953 1197 111 1153 DFRRQJI3VX1 $T=371280 194880 1 180 $X=355730 $Y=194240
X8980 3 1 161 170 105 1291 DFRRQJI3VX1 $T=363440 78400 1 0 $X=363010 $Y=73280
X8981 3 1 161 169 105 741 DFRRQJI3VX1 $T=378560 78400 1 180 $X=363010 $Y=77760
X8982 3 1 161 739 105 1293 DFRRQJI3VX1 $T=363440 87360 0 0 $X=363010 $Y=86720
X8983 3 1 161 754 105 956 DFRRQJI3VX1 $T=363440 96320 1 0 $X=363010 $Y=91200
X8984 3 1 161 756 111 734 DFRRQJI3VX1 $T=378560 150080 1 180 $X=363010 $Y=149440
X8985 3 1 161 755 111 1292 DFRRQJI3VX1 $T=363440 159040 1 0 $X=363010 $Y=153920
X8986 3 1 154 757 105 165 DFRRQJI3VX1 $T=379120 42560 0 180 $X=363570 $Y=37440
X8987 3 1 154 758 105 1288 DFRRQJI3VX1 $T=379120 42560 1 180 $X=363570 $Y=41920
X8988 3 1 154 748 105 164 DFRRQJI3VX1 $T=379120 51520 0 180 $X=363570 $Y=46400
X8989 3 1 154 749 105 730 DFRRQJI3VX1 $T=379120 60480 0 180 $X=363570 $Y=55360
X8990 3 1 154 752 105 955 DFRRQJI3VX1 $T=364000 69440 0 0 $X=363570 $Y=68800
X8991 3 1 161 745 111 1158 DFRRQJI3VX1 $T=364000 159040 0 0 $X=363570 $Y=158400
X8992 3 1 161 759 111 1155 DFRRQJI3VX1 $T=379120 168000 0 180 $X=363570 $Y=162880
X8993 3 1 161 750 111 1154 DFRRQJI3VX1 $T=379120 168000 1 180 $X=363570 $Y=167360
X8994 3 1 154 751 105 1412 DFRRQJI3VX1 $T=379680 33600 1 180 $X=364130 $Y=32960
X8995 3 1 154 753 105 174 DFRRQJI3VX1 $T=367360 69440 1 0 $X=366930 $Y=64320
X8996 3 1 772 1413 1208 210 957 ON211JI3VX1 $T=53200 69440 0 180 $X=48850 $Y=64320
X8997 3 1 16 1211 774 209 222 ON211JI3VX1 $T=52080 51520 0 0 $X=51650 $Y=50880
X8998 3 1 222 997 7 210 enable ON211JI3VX1 $T=54320 60480 0 0 $X=53890 $Y=59840
X8999 3 1 242 999 1003 998 781 ON211JI3VX1 $T=58800 185920 0 180 $X=54450 $Y=180800
X9000 3 1 35 1000 1392 784 780 ON211JI3VX1 $T=60480 96320 0 180 $X=56130 $Y=91200
X9001 3 1 35 19 1366 788 1006 ON211JI3VX1 $T=65520 96320 0 180 $X=61170 $Y=91200
X9002 3 1 236 1299 1414 790 239 ON211JI3VX1 $T=62160 185920 1 0 $X=61730 $Y=180800
X9003 3 1 35 1012 233 792 791 ON211JI3VX1 $T=71120 96320 0 180 $X=66770 $Y=91200
X9004 3 1 242 1218 1023 250 1020 ON211JI3VX1 $T=75040 185920 0 0 $X=74610 $Y=185280
X9005 3 1 1027 279 1415 259 807 ON211JI3VX1 $T=80080 176960 0 0 $X=79650 $Y=176320
X9006 3 1 enable 1416 312 823 35 ON211JI3VX1 $T=105280 176960 1 180 $X=100930 $Y=176320
X9007 3 1 403 1375 1057 409 1303 ON211JI3VX1 $T=151200 185920 1 180 $X=146850 $Y=185280
X9008 3 1 965 1311 1417 484 876 ON211JI3VX1 $T=204400 194880 1 180 $X=200050 $Y=194240
X9009 3 1 1128 138 658 917 132 ON211JI3VX1 $T=301840 176960 1 0 $X=301410 $Y=171840
X9010 3 1 718 933 1391 1325 696 ON211JI3VX1 $T=331520 176960 1 0 $X=331090 $Y=171840
X9011 3 1 153 689 1143 930 enable ON211JI3VX1 $T=335440 185920 0 180 $X=331090 $Y=180800
X9012 3 1 982 7 976 6 186 ON22JI3VX1 $T=34720 69440 1 180 $X=29810 $Y=68800
X9013 3 1 55 18 1160 777 244 ON22JI3VX1 $T=57120 42560 0 180 $X=52210 $Y=37440
X9014 3 1 232 1013 1418 803 1007 ON22JI3VX1 $T=69440 203840 1 180 $X=64530 $Y=203200
X9015 3 1 1055 355 1419 846 840 ON22JI3VX1 $T=140560 185920 1 0 $X=140130 $Y=180800
X9016 3 1 848 60 1343 847 846 ON22JI3VX1 $T=148960 203840 1 180 $X=144050 $Y=203200
X9017 3 1 855 60 1347 1344 1064 ON22JI3VX1 $T=156800 203840 0 0 $X=156370 $Y=203200
X9018 3 1 963 60 1348 868 1075 ON22JI3VX1 $T=179760 203840 0 180 $X=174850 $Y=198720
X9019 3 1 473 94 1370 489 77 ON22JI3VX1 $T=189280 203840 1 0 $X=188850 $Y=198720
X9020 3 1 473 1237 483 77 474 ON22JI3VX1 $T=193760 203840 1 0 $X=193330 $Y=198720
X9021 3 1 885 506 1350 100 507 ON22JI3VX1 $T=220080 194880 0 0 $X=219650 $Y=194240
X9022 3 1 520 1094 537 890 103 ON22JI3VX1 $T=229600 203840 0 0 $X=229170 $Y=203200
X9023 3 1 553 1420 892 895 894 ON22JI3VX1 $T=246400 194880 0 180 $X=241490 $Y=189760
X9024 3 1 1125 1126 1358 678 920 ON22JI3VX1 $T=304640 194880 1 0 $X=304210 $Y=189760
X9025 3 1 142 139 925 698 665 ON22JI3VX1 $T=316960 185920 1 180 $X=312050 $Y=185280
X9026 3 1 931 928 1137 688 152 ON22JI3VX1 $T=324800 185920 1 0 $X=324370 $Y=180800
X9027 3 1 727 706 1373 940 1153 ON22JI3VX1 $T=347200 194880 1 0 $X=346770 $Y=189760
X9028 3 1 1155 971 729 1330 1154 ON22JI3VX1 $T=361200 176960 0 180 $X=356290 $Y=171840
X9029 3 1 161 1290 111 951 DFRRQJI3VX2 $T=372400 194880 0 180 $X=355730 $Y=189760
X9030 3 1 326 8 192 183 EO3JI3VX1 $T=49840 105280 0 180 $X=38770 $Y=100160
X9031 3 1 326 11 1205 1159 EO3JI3VX1 $T=53760 105280 1 180 $X=42690 $Y=104640
X9032 3 1 985 766 18 NO2JI3VX0 $T=44800 51520 0 180 $X=42130 $Y=46400
X9033 3 1 1421 985 997 NO2JI3VX0 $T=43120 60480 0 0 $X=42690 $Y=59840
X9034 3 1 768 194 196 NO2JI3VX0 $T=43120 78400 1 0 $X=42690 $Y=73280
X9035 3 1 777 993 10 NO2JI3VX0 $T=52640 42560 0 180 $X=49970 $Y=37440
X9036 3 1 1422 1208 16 NO2JI3VX0 $T=51520 60480 1 0 $X=51090 $Y=55360
X9037 3 1 199 958 261 NO2JI3VX0 $T=51520 203840 1 0 $X=51090 $Y=198720
X9038 3 1 778 777 18 NO2JI3VX0 $T=52640 42560 0 0 $X=52210 $Y=41920
X9039 3 1 218 1003 1004 NO2JI3VX0 $T=61040 176960 1 180 $X=58370 $Y=176320
X9040 3 1 231 1161 1015 NO2JI3VX0 $T=68320 194880 1 0 $X=67890 $Y=189760
X9041 3 1 796 1415 236 NO2JI3VX0 $T=71680 176960 0 0 $X=71250 $Y=176320
X9042 3 1 800 25 206 NO2JI3VX0 $T=76720 212800 0 180 $X=74050 $Y=207680
X9043 3 1 286 800 247 NO2JI3VX0 $T=80080 212800 0 180 $X=77410 $Y=207680
X9044 3 1 1040 284 818 NO2JI3VX0 $T=95200 114240 0 180 $X=92530 $Y=109120
X9045 3 1 46 49 48 NO2JI3VX0 $T=113120 194880 1 0 $X=112690 $Y=189760
X9046 3 1 308 1368 38 NO2JI3VX0 $T=113120 194880 0 0 $X=112690 $Y=194240
X9047 3 1 246 451 48 NO2JI3VX0 $T=131600 194880 1 180 $X=128930 $Y=194240
X9048 3 1 1229 388 394 NO2JI3VX0 $T=151760 194880 1 180 $X=149090 $Y=194240
X9049 3 1 394 851 854 NO2JI3VX0 $T=150640 194880 1 0 $X=150210 $Y=189760
X9050 3 1 1064 387 1063 NO2JI3VX0 $T=160720 185920 0 180 $X=158050 $Y=180800
X9051 3 1 63 59 420 NO2JI3VX0 $T=164080 194880 1 180 $X=161410 $Y=194240
X9052 3 1 448 866 1074 NO2JI3VX0 $T=175840 185920 1 180 $X=173170 $Y=185280
X9053 3 1 448 452 75 NO2JI3VX0 $T=185920 203840 0 180 $X=183250 $Y=198720
X9054 3 1 878 1313 509 NO2JI3VX0 $T=210560 194880 0 180 $X=207890 $Y=189760
X9055 3 1 506 1239 99 NO2JI3VX0 $T=224560 194880 0 0 $X=224130 $Y=194240
X9056 3 1 570 1423 1102 NO2JI3VX0 $T=246400 24640 0 0 $X=245970 $Y=24000
X9057 3 1 1249 1105 966 NO2JI3VX0 $T=250880 24640 0 0 $X=250450 $Y=24000
X9058 3 1 575 1107 567 NO2JI3VX0 $T=260960 33600 0 180 $X=258290 $Y=28480
X9059 3 1 104 1424 571 NO2JI3VX0 $T=263200 24640 1 180 $X=260530 $Y=24000
X9060 3 1 620 627 1120 NO2JI3VX0 $T=283360 212800 1 0 $X=282930 $Y=207680
X9061 3 1 1321 1357 627 NO2JI3VX0 $T=291760 212800 1 0 $X=291330 $Y=207680
X9062 3 1 1123 1126 48 NO2JI3VX0 $T=297360 194880 0 0 $X=296930 $Y=194240
X9063 3 1 678 1123 912 NO2JI3VX0 $T=302960 194880 1 180 $X=300290 $Y=194240
X9064 3 1 134 1131 916 NO2JI3VX0 $T=309680 185920 0 180 $X=307010 $Y=180800
X9065 3 1 658 667 134 NO2JI3VX0 $T=310800 185920 1 180 $X=308130 $Y=185280
X9066 3 1 924 1425 138 NO2JI3VX0 $T=313600 176960 0 0 $X=313170 $Y=176320
X9067 3 1 698 1149 139 NO2JI3VX0 $T=335440 185920 1 0 $X=335010 $Y=180800
X9068 3 1 1146 1144 713 NO2JI3VX0 $T=337680 185920 1 180 $X=335010 $Y=185280
X9069 3 1 139 162 1274 NO2JI3VX0 $T=338800 168000 1 180 $X=336130 $Y=167360
X9070 3 1 706 690 714 NO2JI3VX0 $T=343280 185920 0 180 $X=340610 $Y=180800
X9071 3 1 943 939 944 NO2JI3VX0 $T=347760 176960 0 180 $X=345090 $Y=171840
X9072 3 1 1408 6 974 981 ON21JI3VX1 $T=34720 60480 0 0 $X=34290 $Y=59840
X9073 3 1 186 194 983 982 ON21JI3VX1 $T=35840 69440 0 0 $X=35410 $Y=68800
X9074 3 1 1386 200 977 980 ON21JI3VX1 $T=40320 203840 1 180 $X=36530 $Y=203200
X9075 3 1 979 194 764 1203 ON21JI3VX1 $T=44800 69440 0 180 $X=41010 $Y=64320
X9076 3 1 1409 213 1204 990 ON21JI3VX1 $T=46480 33600 1 180 $X=42690 $Y=32960
X9077 3 1 993 1160 990 13 ON21JI3VX1 $T=51520 33600 1 180 $X=47730 $Y=32960
X9078 3 1 218 208 781 1004 ON21JI3VX1 $T=54320 176960 0 0 $X=53890 $Y=176320
X9079 3 1 958 1210 786 1297 ON21JI3VX1 $T=54320 194880 0 0 $X=53890 $Y=194240
X9080 3 1 244 213 789 1362 ON21JI3VX1 $T=61600 33600 0 0 $X=61170 $Y=32960
X9081 3 1 796 25 1018 959 ON21JI3VX1 $T=70560 203840 1 0 $X=70130 $Y=198720
X9082 3 1 1387 286 830 1337 ON21JI3VX1 $T=100240 212800 0 0 $X=99810 $Y=212160
X9083 3 1 107 1046 589 1374 ON21JI3VX1 $T=101920 24640 1 0 $X=101490 $Y=19520
X9084 3 1 829 294 1340 828 ON21JI3VX1 $T=105280 194880 1 180 $X=101490 $Y=194240
X9085 3 1 314 313 1341 312 ON21JI3VX1 $T=122080 185920 1 180 $X=118290 $Y=185280
X9086 3 1 1388 60 1051 1052 ON21JI3VX1 $T=132160 203840 1 180 $X=128370 $Y=203200
X9087 3 1 107 1426 904 1226 ON21JI3VX1 $T=129920 24640 0 0 $X=129490 $Y=24000
X9088 3 1 107 1427 612 841 ON21JI3VX1 $T=141120 33600 1 0 $X=140690 $Y=28480
X9089 3 1 107 1428 602 400 ON21JI3VX1 $T=154000 33600 0 0 $X=153570 $Y=32960
X9090 3 1 413 866 1429 424 ON21JI3VX1 $T=171920 194880 0 180 $X=168130 $Y=189760
X9091 3 1 448 868 436 1234 ON21JI3VX1 $T=171360 203840 1 0 $X=170930 $Y=198720
X9092 3 1 872 77 1236 477 ON21JI3VX1 $T=194320 194880 1 0 $X=193890 $Y=189760
X9093 3 1 107 1085 567 879 ON21JI3VX1 $T=201040 33600 1 0 $X=200610 $Y=28480
X9094 3 1 482 1389 1351 493 ON21JI3VX1 $T=207760 185920 0 0 $X=207330 $Y=185280
X9095 3 1 107 1430 571 1314 ON21JI3VX1 $T=221760 24640 0 0 $X=221330 $Y=24000
X9096 3 1 107 888 575 1241 ON21JI3VX1 $T=226240 33600 1 0 $X=225810 $Y=28480
X9097 3 1 516 1390 1177 1353 ON21JI3VX1 $T=227360 194880 1 0 $X=226930 $Y=189760
X9098 3 1 520 94 1246 890 ON21JI3VX1 $T=229600 203840 1 0 $X=229170 $Y=198720
X9099 3 1 107 1099 104 1245 ON21JI3VX1 $T=236320 33600 0 0 $X=235890 $Y=32960
X9100 3 1 107 1431 1249 1354 ON21JI3VX1 $T=239120 24640 1 0 $X=238690 $Y=19520
X9101 3 1 86 1246 1432 1315 ON21JI3VX1 $T=240800 203840 1 0 $X=240370 $Y=198720
X9102 3 1 107 1433 1102 1355 ON21JI3VX1 $T=247520 42560 0 180 $X=243730 $Y=37440
X9103 3 1 107 1317 966 1316 ON21JI3VX1 $T=256480 33600 1 180 $X=252690 $Y=32960
X9104 3 1 107 1108 570 1110 ON21JI3VX1 $T=258160 33600 0 0 $X=257730 $Y=32960
X9105 3 1 134 1126 1129 1266 ON21JI3VX1 $T=308000 194880 1 180 $X=304210 $Y=194240
X9106 3 1 1131 676 1377 654 ON21JI3VX1 $T=311360 176960 1 180 $X=307570 $Y=176320
X9107 3 1 678 1270 1275 1271 ON21JI3VX1 $T=329280 203840 0 0 $X=328850 $Y=203200
X9108 3 1 612 1065 1434 632 602 OR4JI3VX1 $T=286160 24640 1 180 $X=279570 $Y=24000
X9109 3 1 150 137 1269 663 650 OR4JI3VX1 $T=315840 33600 0 180 $X=309250 $Y=28480
X9110 3 1 704 1139 660 680 478 OR4JI3VX1 $T=331520 24640 1 180 $X=324930 $Y=24000
X9111 3 1 719 947 948 736 946 OR4JI3VX1 $T=353360 33600 0 180 $X=346770 $Y=28480
X9112 3 1 480 494 BUJI3VX16 $T=183120 221760 1 0 $X=182690 $Y=216640
X9113 3 1 131 161 BUJI3VX16 $T=332640 221760 0 180 $X=315970 $Y=216640
X9114 3 1 984 107 BUJI3VX6 $T=37520 78400 1 180 $X=30370 $Y=77760
X9115 3 1 131 1267 BUJI3VX6 $T=309680 221760 1 0 $X=309250 $Y=216640
X9116 3 1 979 7 6 1364 1435 ON31JI3VX1 $T=35840 69440 0 180 $X=30930 $Y=64320
X9117 3 1 10 209 213 190 1436 ON31JI3VX1 $T=47040 42560 0 180 $X=42130 $Y=37440
X9118 3 1 199 992 200 1335 1296 ON31JI3VX1 $T=52080 203840 1 180 $X=47170 $Y=203200
X9119 3 1 282 281 286 1032 1437 ON31JI3VX1 $T=90160 212800 0 180 $X=85250 $Y=207680
X9120 3 1 369 843 60 360 1054 ON31JI3VX1 $T=144480 203840 1 180 $X=139570 $Y=203200
X9121 3 1 852 1229 60 844 1058 ON31JI3VX1 $T=152880 212800 0 180 $X=147970 $Y=207680
X9122 3 1 426 63 60 1066 1345 ON31JI3VX1 $T=166320 203840 1 180 $X=161410 $Y=203200
X9123 3 1 885 498 94 1349 1091 ON31JI3VX1 $T=223440 203840 1 180 $X=218530 $Y=203200
X9124 3 1 522 103 1094 546 1371 ON31JI3VX1 $T=231840 194880 0 0 $X=231410 $Y=194240
X9125 3 1 142 926 678 679 1324 ON31JI3VX1 $T=329280 203840 1 180 $X=324370 $Y=203200
X9126 3 1 701 678 1141 1276 970 ON31JI3VX1 $T=332640 203840 0 0 $X=332210 $Y=203200
X9127 3 1 727 942 678 1200 1281 ON31JI3VX1 $T=344400 203840 1 0 $X=343970 $Y=198720
X9128 3 1 551 535 DLY4JI3VX1 $T=232960 212800 0 0 $X=232530 $Y=212160
X9129 3 1 SPI_CS 581 DLY4JI3VX1 $T=258720 221760 1 0 $X=258290 $Y=216640
X9130 3 1 55 76 107 NO2I1JI3VX2 $T=192640 42560 0 180 $X=187170 $Y=37440
X9131 3 1 131 604 BUJI3VX12 $T=275520 150080 1 0 $X=275090 $Y=144960
X9132 3 1 131 633 BUJI3VX12 $T=287840 150080 1 0 $X=287410 $Y=144960
X9133 3 1 609 up_switches<22> INJI3VX3 $T=281680 24640 1 0 $X=281250 $Y=19520
X9134 3 1 649 404 INJI3VX3 $T=304080 42560 1 0 $X=303650 $Y=37440
X9135 3 1 740 up_switches<3> INJI3VX3 $T=367360 24640 1 0 $X=366930 $Y=19520
X9136 3 1 746 up_switches<2> INJI3VX3 $T=370720 24640 1 0 $X=370290 $Y=19520
X9137 3 1 1438 1421 772 991 957 NA4JI3VX0 $T=50400 60480 1 180 $X=46050 $Y=59840
X9138 3 1 828 1339 447 829 1439 NA4JI3VX0 $T=100800 185920 0 0 $X=100370 $Y=185280
X9139 3 1 1423 1180 1424 1107 1105 NA4JI3VX0 $T=255360 24640 0 0 $X=254930 $Y=24000
X9140 3 1 609 1187 746 740 625 NA4JI3VX0 $T=288960 24640 0 0 $X=288530 $Y=24000
X9141 3 1 929 464 1136 1360 1425 NA4JI3VX0 $T=329280 176960 1 180 $X=324930 $Y=176320
X9142 3 1 1213 1299 1393 294 OR3JI3VX1 $T=63840 194880 1 0 $X=63410 $Y=189760
X9143 3 1 589 904 644 1116 OR3JI3VX1 $T=272720 24640 1 0 $X=272290 $Y=19520
X9144 3 1 948 1152 1284 673 OR3JI3VX1 $T=349440 24640 1 180 $X=345090 $Y=24000
X9145 3 1 1116 625 1434 1180 NO3JI3VX1 $T=274960 24640 0 0 $X=274530 $Y=24000
X9146 3 1 973 1333 179 379 216 FAJI3VX1 $T=23520 132160 0 0 $X=23090 $Y=131520
X9147 3 1 972 978 5 345 1333 FAJI3VX1 $T=23520 150080 0 0 $X=23090 $Y=149440
X9148 3 1 975 1365 204 331 192 FAJI3VX1 $T=25200 105280 0 0 $X=24770 $Y=104640
X9149 3 1 760 1021 182 986 1365 FAJI3VX1 $T=25200 114240 1 0 $X=24770 $Y=109120
X9150 3 1 779 987 197 345 770 FAJI3VX1 $T=53760 150080 1 180 $X=38770 $Y=149440
X9151 3 1 1212 770 198 379 219 FAJI3VX1 $T=54320 150080 0 180 $X=39330 $Y=144960
X9152 3 1 15 775 20 331 1205 FAJI3VX1 $T=40880 114240 1 0 $X=40450 $Y=109120
X9153 3 1 17 229 782 986 775 FAJI3VX1 $T=40880 114240 0 0 $X=40450 $Y=113600
X9154 3 1 233 211 204 1440 996 FAJI3VX1 $T=41440 96320 0 0 $X=41010 $Y=95680
X9155 3 1 1366 1336 182 205 211 FAJI3VX1 $T=65520 105280 0 180 $X=50530 $Y=100160
X9156 3 1 1001 216 795 373 240 FAJI3VX1 $T=56560 132160 0 0 $X=56130 $Y=131520
X9157 3 1 23 254 793 333 229 FAJI3VX1 $T=58240 114240 0 0 $X=57810 $Y=113600
X9158 3 1 1002 219 237 373 21 FAJI3VX1 $T=58240 150080 1 0 $X=57810 $Y=144960
X9159 3 1 249 806 256 333 1021 FAJI3VX1 $T=68320 105280 0 0 $X=67890 $Y=104640
X9160 3 1 798 240 263 842 1025 FAJI3VX1 $T=70560 132160 1 0 $X=70130 $Y=127040
X9161 3 1 799 21 31 842 1026 FAJI3VX1 $T=70560 141120 1 0 $X=70130 $Y=136000
X9162 3 1 801 1026 26 1037 254 FAJI3VX1 $T=72800 123200 1 0 $X=72370 $Y=118080
X9163 3 1 1022 1025 270 1037 806 FAJI3VX1 $T=74480 114240 0 0 $X=74050 $Y=113600
X9164 3 1 891 116 BUJI3VX4 $T=233520 114240 0 180 $X=227490 $Y=109120
X9165 3 1 1305 434 INJI3VX1 $T=170800 185920 1 0 $X=170370 $Y=180800
X9166 3 1 503 499 INJI3VX1 $T=223440 221760 0 180 $X=221330 $Y=216640
X9167 3 1 499 185 DLY2JI3VX1 $T=175840 221760 1 0 $X=175410 $Y=216640
X9168 3 1 565 126 DLY2JI3VX1 $T=256480 212800 0 0 $X=256050 $Y=212160
X9169 3 1 208 195 185 24 4 208 SDFRRQJI3VX1 $T=42560 176960 1 180 $X=21970 $Y=176320
X9170 3 1 766 18 180 985 14 18 SDFRRQJI3VX1 $T=43120 42560 1 180 $X=22530 $Y=41920
X9171 3 1 44 28 180 41 322 28 SDFRRQJI3VX1 $T=101360 60480 0 180 $X=80770 $Y=55360
X9172 3 1 44 289 180 343 322 289 SDFRRQJI3VX1 $T=101360 60480 1 180 $X=80770 $Y=59840
X9173 3 1 307 41 180 251 322 251 SDFRRQJI3VX1 $T=101360 69440 0 180 $X=80770 $Y=64320
X9174 3 1 307 40 180 287 322 287 SDFRRQJI3VX1 $T=101360 69440 1 180 $X=80770 $Y=68800
X9175 3 1 307 343 180 288 322 288 SDFRRQJI3VX1 $T=101360 78400 0 180 $X=80770 $Y=73280
X9176 3 1 43 295 180 343 322 295 SDFRRQJI3VX1 $T=105280 51520 1 180 $X=84690 $Y=50880
X9177 3 1 45 297 180 41 322 297 SDFRRQJI3VX1 $T=105280 132160 0 180 $X=84690 $Y=127040
X9178 3 1 45 298 180 343 322 298 SDFRRQJI3VX1 $T=105280 132160 1 180 $X=84690 $Y=131520
X9179 3 1 45 299 180 40 322 299 SDFRRQJI3VX1 $T=105280 141120 0 180 $X=84690 $Y=136000
X9180 3 1 45 30 180 303 322 30 SDFRRQJI3VX1 $T=105280 141120 1 180 $X=84690 $Y=140480
X9181 3 1 43 340 53 41 322 340 SDFRRQJI3VX1 $T=113120 60480 1 0 $X=112690 $Y=55360
X9182 3 1 43 341 53 40 322 341 SDFRRQJI3VX1 $T=113120 60480 0 0 $X=112690 $Y=59840
X9183 3 1 44 306 53 40 322 306 SDFRRQJI3VX1 $T=113120 69440 1 0 $X=112690 $Y=64320
X9184 3 1 44 352 56 336 322 352 SDFRRQJI3VX1 $T=113120 69440 0 0 $X=112690 $Y=68800
X9185 3 1 44 342 53 303 322 342 SDFRRQJI3VX1 $T=113120 87360 1 0 $X=112690 $Y=82240
X9186 3 1 322 40 53 343 116 40 SDFRRQJI3VX1 $T=113120 114240 0 0 $X=112690 $Y=113600
X9187 3 1 322 41 53 40 116 41 SDFRRQJI3VX1 $T=113120 123200 0 0 $X=112690 $Y=122560
X9188 3 1 322 343 53 303 116 343 SDFRRQJI3VX1 $T=113120 132160 1 0 $X=112690 $Y=127040
X9189 3 1 322 303 53 336 116 303 SDFRRQJI3VX1 $T=113120 132160 0 0 $X=112690 $Y=131520
X9190 3 1 322 336 53 397 116 336 SDFRRQJI3VX1 $T=113120 141120 1 0 $X=112690 $Y=136000
X9191 3 1 307 303 53 339 322 339 SDFRRQJI3VX1 $T=113120 141120 0 0 $X=112690 $Y=140480
X9192 3 1 45 344 53 397 322 344 SDFRRQJI3VX1 $T=113120 150080 1 0 $X=112690 $Y=144960
X9193 3 1 45 304 53 336 322 304 SDFRRQJI3VX1 $T=113120 159040 1 0 $X=112690 $Y=153920
X9194 3 1 307 336 53 349 322 349 SDFRRQJI3VX1 $T=115920 159040 0 0 $X=115490 $Y=158400
X9195 3 1 43 358 53 303 322 358 SDFRRQJI3VX1 $T=120960 78400 0 0 $X=120530 $Y=77760
X9196 3 1 43 375 56 336 322 375 SDFRRQJI3VX1 $T=125440 78400 1 0 $X=125010 $Y=73280
X9197 3 1 45 364 56 65 322 364 SDFRRQJI3VX1 $T=145600 96320 1 180 $X=125010 $Y=95680
X9198 3 1 307 397 53 337 322 337 SDFRRQJI3VX1 $T=125440 150080 0 0 $X=125010 $Y=149440
X9199 3 1 45 378 53 393 322 378 SDFRRQJI3VX1 $T=148400 96320 0 180 $X=127810 $Y=91200
X9200 3 1 307 65 56 390 322 390 SDFRRQJI3VX1 $T=153440 141120 1 180 $X=132850 $Y=140480
X9201 3 1 307 393 56 391 322 391 SDFRRQJI3VX1 $T=153440 150080 0 180 $X=132850 $Y=144960
X9202 3 1 322 393 53 65 116 393 SDFRRQJI3VX1 $T=133840 123200 0 0 $X=133410 $Y=122560
X9203 3 1 322 397 56 393 116 397 SDFRRQJI3VX1 $T=156240 132160 0 180 $X=135650 $Y=127040
X9204 3 1 43 414 56 393 322 414 SDFRRQJI3VX1 $T=142800 69440 0 0 $X=142370 $Y=68800
X9205 3 1 44 415 56 397 322 415 SDFRRQJI3VX1 $T=142800 87360 1 0 $X=142370 $Y=82240
X9206 3 1 43 418 56 397 322 418 SDFRRQJI3VX1 $T=145040 87360 0 0 $X=144610 $Y=86720
X9207 3 1 44 396 56 393 322 396 SDFRRQJI3VX1 $T=147280 78400 1 0 $X=146850 $Y=73280
X9208 3 1 45 370 56 433 322 370 SDFRRQJI3VX1 $T=167440 105280 0 180 $X=146850 $Y=100160
X9209 3 1 45 380 56 72 322 380 SDFRRQJI3VX1 $T=168560 96320 1 180 $X=147970 $Y=95680
X9210 3 1 307 72 56 401 322 401 SDFRRQJI3VX1 $T=175840 141120 1 180 $X=155250 $Y=140480
X9211 3 1 45 1060 56 62 322 1060 SDFRRQJI3VX1 $T=179200 114240 0 180 $X=158610 $Y=109120
X9212 3 1 322 70 71 62 116 70 SDFRRQJI3VX1 $T=159040 132160 1 0 $X=158610 $Y=127040
X9213 3 1 45 406 56 70 322 406 SDFRRQJI3VX1 $T=180320 105280 1 180 $X=159730 $Y=104640
X9214 3 1 322 433 71 70 116 433 SDFRRQJI3VX1 $T=160160 114240 0 0 $X=159730 $Y=113600
X9215 3 1 322 500 71 41 116 500 SDFRRQJI3VX1 $T=160160 123200 0 0 $X=159730 $Y=122560
X9216 3 1 126 72 56 433 116 72 SDFRRQJI3VX1 $T=180880 132160 1 180 $X=160290 $Y=131520
X9217 3 1 322 65 56 72 116 65 SDFRRQJI3VX1 $T=181440 141120 0 180 $X=160850 $Y=136000
X9218 3 1 307 433 56 438 SPI_CS 438 SDFRRQJI3VX1 $T=182000 150080 0 180 $X=161410 $Y=144960
X9219 3 1 307 70 71 449 SPI_CS 449 SDFRRQJI3VX1 $T=164080 150080 0 0 $X=163650 $Y=149440
X9220 3 1 43 454 71 65 SPI_CS 454 SDFRRQJI3VX1 $T=165200 78400 0 0 $X=164770 $Y=77760
X9221 3 1 44 455 71 65 SPI_CS 455 SDFRRQJI3VX1 $T=165760 87360 0 0 $X=165330 $Y=86720
X9222 3 1 44 456 71 72 SPI_CS 456 SDFRRQJI3VX1 $T=165760 96320 1 0 $X=165330 $Y=91200
X9223 3 1 43 67 71 72 SPI_CS 67 SDFRRQJI3VX1 $T=169680 123200 1 0 $X=169250 $Y=118080
X9224 3 1 307 62 71 441 SPI_CS 441 SDFRRQJI3VX1 $T=169680 159040 1 0 $X=169250 $Y=153920
X9225 3 1 43 463 71 433 SPI_CS 463 SDFRRQJI3VX1 $T=171360 96320 0 0 $X=170930 $Y=95680
X9226 3 1 44 1174 71 433 SPI_CS 1174 SDFRRQJI3VX1 $T=171360 105280 1 0 $X=170930 $Y=100160
X9227 3 1 43 1175 71 70 SPI_CS 1175 SDFRRQJI3VX1 $T=185920 87360 0 0 $X=185490 $Y=86720
X9228 3 1 45 458 71 497 SPI_CS 458 SDFRRQJI3VX1 $T=207200 150080 1 180 $X=186610 $Y=149440
X9229 3 1 44 479 71 70 SPI_CS 479 SDFRRQJI3VX1 $T=187600 96320 1 0 $X=187170 $Y=91200
X9230 3 1 43 84 71 500 SPI_CS 84 SDFRRQJI3VX1 $T=208320 105280 1 180 $X=187730 $Y=104640
X9231 3 1 44 87 71 500 SPI_CS 87 SDFRRQJI3VX1 $T=210000 123200 0 180 $X=189410 $Y=118080
X9232 3 1 307 127 71 74 SPI_CS 74 SDFRRQJI3VX1 $T=210000 159040 0 180 $X=189410 $Y=153920
X9233 3 1 45 481 71 500 SPI_CS 481 SDFRRQJI3VX1 $T=211120 132160 0 180 $X=190530 $Y=127040
X9234 3 1 43 95 518 528 SPI_CS 95 SDFRRQJI3VX1 $T=218960 87360 0 0 $X=218530 $Y=86720
X9235 3 1 44 525 518 528 SPI_CS 525 SDFRRQJI3VX1 $T=218960 96320 1 0 $X=218530 $Y=91200
X9236 3 1 43 526 518 497 SPI_CS 526 SDFRRQJI3VX1 $T=218960 96320 0 0 $X=218530 $Y=95680
X9237 3 1 44 96 518 497 SPI_CS 96 SDFRRQJI3VX1 $T=218960 105280 0 0 $X=218530 $Y=104640
X9238 3 1 307 159 536 527 SPI_CS 527 SDFRRQJI3VX1 $T=218960 114240 0 0 $X=218530 $Y=113600
X9239 3 1 126 528 518 497 116 528 SDFRRQJI3VX1 $T=218960 123200 1 0 $X=218530 $Y=118080
X9240 3 1 126 497 518 500 116 497 SDFRRQJI3VX1 $T=218960 123200 0 0 $X=218530 $Y=122560
X9241 3 1 126 62 518 504 116 62 SDFRRQJI3VX1 $T=218960 132160 1 0 $X=218530 $Y=127040
X9242 3 1 126 1100 518 528 116 1100 SDFRRQJI3VX1 $T=218960 132160 0 0 $X=218530 $Y=131520
X9243 3 1 307 605 518 501 SPI_CS 501 SDFRRQJI3VX1 $T=218960 141120 0 0 $X=218530 $Y=140480
X9244 3 1 307 574 518 502 SPI_CS 502 SDFRRQJI3VX1 $T=218960 150080 1 0 $X=218530 $Y=144960
X9245 3 1 45 524 518 1100 SPI_CS 524 SDFRRQJI3VX1 $T=218960 150080 0 0 $X=218530 $Y=149440
X9246 3 1 45 88 518 528 SPI_CS 88 SDFRRQJI3VX1 $T=218960 159040 1 0 $X=218530 $Y=153920
X9247 3 1 307 504 518 529 SPI_CS 529 SDFRRQJI3VX1 $T=218960 159040 0 0 $X=218530 $Y=158400
X9248 3 1 307 608 518 538 SPI_CS 538 SDFRRQJI3VX1 $T=246960 141120 0 180 $X=226370 $Y=136000
X9249 3 1 581 127 108 535 116 127 SDFRRQJI3VX1 $T=227360 221760 1 0 $X=226930 $Y=216640
X9250 3 1 44 102 518 545 SPI_CS 102 SDFRRQJI3VX1 $T=252000 105280 0 180 $X=231410 $Y=100160
X9251 3 1 307 623 518 521 SPI_CS 521 SDFRRQJI3VX1 $T=233520 114240 1 0 $X=233090 $Y=109120
X9252 3 1 45 552 518 545 SPI_CS 552 SDFRRQJI3VX1 $T=253680 168000 0 180 $X=233090 $Y=162880
X9253 3 1 43 568 518 1100 SPI_CS 568 SDFRRQJI3VX1 $T=239120 87360 0 0 $X=238690 $Y=86720
X9254 3 1 44 569 518 1100 SPI_CS 569 SDFRRQJI3VX1 $T=239120 96320 1 0 $X=238690 $Y=91200
X9255 3 1 45 893 536 561 SPI_CS 893 SDFRRQJI3VX1 $T=259280 150080 0 180 $X=238690 $Y=144960
X9256 3 1 307 645 518 530 SPI_CS 530 SDFRRQJI3VX1 $T=259280 150080 1 180 $X=238690 $Y=149440
X9257 3 1 45 110 536 566 SPI_CS 110 SDFRRQJI3VX1 $T=259280 159040 0 180 $X=238690 $Y=153920
X9258 3 1 43 572 536 545 SPI_CS 572 SDFRRQJI3VX1 $T=240240 105280 0 0 $X=239810 $Y=104640
X9259 3 1 307 125 518 531 SPI_CS 531 SDFRRQJI3VX1 $T=260400 114240 1 180 $X=239810 $Y=113600
X9260 3 1 307 742 518 532 SPI_CS 532 SDFRRQJI3VX1 $T=260400 123200 0 180 $X=239810 $Y=118080
X9261 3 1 307 684 518 564 SPI_CS 564 SDFRRQJI3VX1 $T=260400 123200 1 180 $X=239810 $Y=122560
X9262 3 1 126 566 108 1100 116 566 SDFRRQJI3VX1 $T=240800 132160 1 0 $X=240370 $Y=127040
X9263 3 1 126 561 108 566 116 561 SDFRRQJI3VX1 $T=261520 132160 1 180 $X=240930 $Y=131520
X9264 3 1 126 545 108 561 116 545 SDFRRQJI3VX1 $T=241920 141120 0 0 $X=241490 $Y=140480
X9265 3 1 126 583 108 1104 116 583 SDFRRQJI3VX1 $T=248080 212800 1 0 $X=247650 $Y=207680
X9266 3 1 44 584 518 566 SPI_CS 584 SDFRRQJI3VX1 $T=248640 87360 1 0 $X=248210 $Y=82240
X9267 3 1 43 585 518 561 SPI_CS 585 SDFRRQJI3VX1 $T=249200 78400 1 0 $X=248770 $Y=73280
X9268 3 1 44 586 518 561 SPI_CS 586 SDFRRQJI3VX1 $T=249200 78400 0 0 $X=248770 $Y=77760
X9269 3 1 43 587 518 566 SPI_CS 587 SDFRRQJI3VX1 $T=249200 96320 0 0 $X=248770 $Y=95680
X9270 3 1 126 1104 108 580 116 1104 SDFRRQJI3VX1 $T=269920 203840 0 180 $X=249330 $Y=198720
X9271 3 1 307 737 518 591 SPI_CS 591 SDFRRQJI3VX1 $T=253680 114240 1 0 $X=253250 $Y=109120
X9272 3 1 172 577 108 592 116 577 SDFRRQJI3VX1 $T=274960 168000 0 180 $X=254370 $Y=162880
X9273 3 1 126 1319 108 598 116 580 SDFRRQJI3VX1 $T=275520 194880 1 180 $X=254930 $Y=194240
X9274 3 1 126 592 108 596 116 592 SDFRRQJI3VX1 $T=276080 159040 1 180 $X=255490 $Y=158400
X9275 3 1 126 900 131 119 116 598 SDFRRQJI3VX1 $T=255920 194880 1 0 $X=255490 $Y=189760
X9276 3 1 126 1250 131 577 116 1114 SDFRRQJI3VX1 $T=257600 168000 0 0 $X=257170 $Y=167360
X9277 3 1 172 1256 108 1114 116 119 SDFRRQJI3VX1 $T=277760 176960 0 180 $X=257170 $Y=171840
X9278 3 1 45 573 536 596 SPI_CS 573 SDFRRQJI3VX1 $T=279440 159040 0 180 $X=258850 $Y=153920
X9279 3 1 43 123 536 596 SPI_CS 123 SDFRRQJI3VX1 $T=284480 105280 1 180 $X=263890 $Y=104640
X9280 3 1 126 742 108 159 116 742 SDFRRQJI3VX1 $T=264320 123200 1 0 $X=263890 $Y=118080
X9281 3 1 126 125 108 737 116 125 SDFRRQJI3VX1 $T=264320 123200 0 0 $X=263890 $Y=122560
X9282 3 1 126 596 108 545 116 596 SDFRRQJI3VX1 $T=264320 141120 1 0 $X=263890 $Y=136000
X9283 3 1 126 684 108 608 116 684 SDFRRQJI3VX1 $T=264880 132160 1 0 $X=264450 $Y=127040
X9284 3 1 172 608 108 574 116 608 SDFRRQJI3VX1 $T=264880 132160 0 0 $X=264450 $Y=131520
X9285 3 1 172 574 108 605 116 574 SDFRRQJI3VX1 $T=285600 141120 1 180 $X=265010 $Y=140480
X9286 3 1 44 615 536 62 172 615 SDFRRQJI3VX1 $T=269920 96320 0 0 $X=269490 $Y=95680
X9287 3 1 43 619 536 62 172 619 SDFRRQJI3VX1 $T=270480 96320 1 0 $X=270050 $Y=91200
X9288 3 1 44 621 154 574 172 621 SDFRRQJI3VX1 $T=272160 87360 1 0 $X=271730 $Y=82240
X9289 3 1 43 622 154 574 172 622 SDFRRQJI3VX1 $T=272160 87360 0 0 $X=271730 $Y=86720
X9290 3 1 45 636 154 574 172 636 SDFRRQJI3VX1 $T=277760 159040 0 0 $X=277330 $Y=158400
X9291 3 1 45 638 154 127 172 638 SDFRRQJI3VX1 $T=279440 159040 1 0 $X=279010 $Y=153920
X9292 3 1 172 737 154 623 116 737 SDFRRQJI3VX1 $T=288400 123200 1 0 $X=287970 $Y=118080
X9293 3 1 172 623 154 742 116 623 SDFRRQJI3VX1 $T=288400 123200 0 0 $X=287970 $Y=122560
X9294 3 1 172 645 154 125 116 645 SDFRRQJI3VX1 $T=288400 132160 1 0 $X=287970 $Y=127040
X9295 3 1 43 651 154 608 172 651 SDFRRQJI3VX1 $T=288960 78400 1 0 $X=288530 $Y=73280
X9296 3 1 43 652 154 127 172 652 SDFRRQJI3VX1 $T=288960 105280 0 0 $X=288530 $Y=104640
X9297 3 1 44 653 154 127 172 653 SDFRRQJI3VX1 $T=288960 114240 1 0 $X=288530 $Y=109120
X9298 3 1 172 159 154 684 116 159 SDFRRQJI3VX1 $T=288960 132160 0 0 $X=288530 $Y=131520
X9299 3 1 172 605 154 127 116 605 SDFRRQJI3VX1 $T=288960 141120 1 0 $X=288530 $Y=136000
X9300 3 1 172 504 154 645 116 504 SDFRRQJI3VX1 $T=309120 141120 1 180 $X=288530 $Y=140480
X9301 3 1 44 656 154 608 172 656 SDFRRQJI3VX1 $T=289520 78400 0 0 $X=289090 $Y=77760
X9302 3 1 45 136 154 608 172 136 SDFRRQJI3VX1 $T=289520 150080 0 0 $X=289090 $Y=149440
X9303 3 1 44 666 536 596 SPI_CS 666 SDFRRQJI3VX1 $T=292320 114240 0 0 $X=291890 $Y=113600
X9304 3 1 44 709 154 504 172 709 SDFRRQJI3VX1 $T=324800 69440 0 0 $X=324370 $Y=68800
X9305 3 1 43 710 154 504 172 710 SDFRRQJI3VX1 $T=324800 78400 1 0 $X=324370 $Y=73280
X9306 3 1 43 711 154 645 172 711 SDFRRQJI3VX1 $T=324800 87360 1 0 $X=324370 $Y=82240
X9307 3 1 44 148 154 645 172 148 SDFRRQJI3VX1 $T=324800 87360 0 0 $X=324370 $Y=86720
X9308 3 1 43 681 154 605 172 681 SDFRRQJI3VX1 $T=324800 114240 0 0 $X=324370 $Y=113600
X9309 3 1 44 683 154 605 172 683 SDFRRQJI3VX1 $T=324800 123200 1 0 $X=324370 $Y=118080
X9310 3 1 43 708 131 684 172 708 SDFRRQJI3VX1 $T=324800 123200 0 0 $X=324370 $Y=122560
X9311 3 1 45 712 154 605 172 712 SDFRRQJI3VX1 $T=324800 132160 1 0 $X=324370 $Y=127040
X9312 3 1 45 149 154 645 172 149 SDFRRQJI3VX1 $T=324800 150080 1 0 $X=324370 $Y=144960
X9313 3 1 45 685 131 504 172 685 SDFRRQJI3VX1 $T=326480 159040 1 0 $X=326050 $Y=153920
X9314 3 1 44 720 131 159 172 720 SDFRRQJI3VX1 $T=336560 114240 1 0 $X=336130 $Y=109120
X9315 3 1 45 721 131 684 172 721 SDFRRQJI3VX1 $T=336560 132160 0 0 $X=336130 $Y=131520
X9316 3 1 45 717 131 159 172 717 SDFRRQJI3VX1 $T=336560 141120 1 0 $X=336130 $Y=136000
X9317 3 1 43 724 131 159 172 724 SDFRRQJI3VX1 $T=337120 105280 0 0 $X=336690 $Y=104640
X9318 3 1 43 728 154 125 172 728 SDFRRQJI3VX1 $T=338240 78400 0 0 $X=337810 $Y=77760
X9319 3 1 44 726 154 125 172 726 SDFRRQJI3VX1 $T=338240 96320 1 0 $X=337810 $Y=91200
X9320 3 1 43 739 131 742 172 739 SDFRRQJI3VX1 $T=344960 123200 1 0 $X=344530 $Y=118080
X9321 3 1 44 1156 131 684 172 1156 SDFRRQJI3VX1 $T=344960 123200 0 0 $X=344530 $Y=122560
X9322 3 1 45 168 131 125 172 168 SDFRRQJI3VX1 $T=344960 132160 1 0 $X=344530 $Y=127040
X9323 3 1 43 752 131 623 172 752 SDFRRQJI3VX1 $T=360640 96320 0 0 $X=360210 $Y=95680
X9324 3 1 44 753 131 623 172 753 SDFRRQJI3VX1 $T=360640 105280 1 0 $X=360210 $Y=100160
X9325 3 1 43 754 131 737 172 754 SDFRRQJI3VX1 $T=360640 114240 1 0 $X=360210 $Y=109120
X9326 3 1 44 170 131 737 172 170 SDFRRQJI3VX1 $T=360640 114240 0 0 $X=360210 $Y=113600
X9327 3 1 45 755 131 623 172 755 SDFRRQJI3VX1 $T=360640 132160 0 0 $X=360210 $Y=131520
X9328 3 1 45 756 131 737 172 756 SDFRRQJI3VX1 $T=360640 141120 1 0 $X=360210 $Y=136000
X9329 3 1 45 745 131 742 172 745 SDFRRQJI3VX1 $T=360640 141120 0 0 $X=360210 $Y=140480
X9330 3 1 44 169 131 742 172 169 SDFRRQJI3VX1 $T=365120 123200 1 0 $X=364690 $Y=118080
X9331 3 1 53 180 BUJI3VX3 $T=100800 168000 1 0 $X=100370 $Y=162880
X9332 3 1 1048 enable BUJI3VX3 $T=122640 185920 0 0 $X=122210 $Y=185280
X9333 3 1 76 649 BUJI3VX3 $T=192640 24640 0 0 $X=192210 $Y=24000
X9334 3 1 131 908 BUJI3VX3 $T=280000 168000 0 0 $X=279570 $Y=167360
X9335 3 1 131 611 BUJI3VX3 $T=280560 168000 1 0 $X=280130 $Y=162880
X9336 3 1 1065 up_switches<18> BUJI3VX3 $T=295680 24640 0 0 $X=295250 $Y=24000
X9337 3 1 131 1261 BUJI3VX3 $T=295680 176960 1 0 $X=295250 $Y=171840
X9338 3 1 632 up_switches<17> BUJI3VX3 $T=299040 24640 1 0 $X=298610 $Y=19520
X9339 3 1 131 913 BUJI3VX3 $T=301280 212800 1 0 $X=300850 $Y=207680
X9340 3 1 644 up_switches<16> BUJI3VX3 $T=302960 24640 1 0 $X=302530 $Y=19520
X9341 3 1 131 659 BUJI3VX3 $T=302960 212800 0 0 $X=302530 $Y=212160
X9342 3 1 131 919 BUJI3VX3 $T=303520 150080 1 0 $X=303090 $Y=144960
X9343 3 1 131 1132 BUJI3VX3 $T=306880 176960 1 0 $X=306450 $Y=171840
X9344 3 1 650 up_switches<15> BUJI3VX3 $T=307440 24640 1 0 $X=307010 $Y=19520
X9345 3 1 663 up_switches<14> BUJI3VX3 $T=311360 24640 1 0 $X=310930 $Y=19520
X9346 3 1 131 677 BUJI3VX3 $T=313600 203840 0 0 $X=313170 $Y=203200
X9347 3 1 478 up_switches<13> BUJI3VX3 $T=327600 24640 0 180 $X=323250 $Y=19520
X9348 3 1 680 up_switches<12> BUJI3VX3 $T=337120 24640 1 180 $X=332770 $Y=24000
X9349 3 1 131 700 BUJI3VX3 $T=334880 159040 0 0 $X=334450 $Y=158400
X9350 3 1 704 up_switches<11> BUJI3VX3 $T=341040 24640 0 180 $X=336690 $Y=19520
X9351 3 1 1139 up_switches<10> BUJI3VX3 $T=341040 24640 1 180 $X=336690 $Y=24000
X9352 3 1 946 up_switches<9> BUJI3VX3 $T=344960 24640 1 180 $X=340610 $Y=24000
X9353 3 1 947 up_switches<8> BUJI3VX3 $T=348880 24640 0 180 $X=344530 $Y=19520
X9354 3 1 1152 up_switches<7> BUJI3VX3 $T=352800 24640 0 180 $X=348450 $Y=19520
X9355 3 1 1284 up_switches<6> BUJI3VX3 $T=352240 24640 0 0 $X=351810 $Y=24000
X9356 3 1 719 up_switches<5> BUJI3VX3 $T=353360 24640 1 0 $X=352930 $Y=19520
X9357 3 1 131 1287 BUJI3VX3 $T=355040 203840 0 0 $X=354610 $Y=203200
X9358 3 1 131 953 BUJI3VX3 $T=358960 203840 0 0 $X=358530 $Y=203200
X9359 3 1 736 up_switches<4> BUJI3VX3 $T=364560 24640 1 180 $X=360210 $Y=24000
X9360 3 1 150 up_switches<1> BUJI3VX3 $T=374080 24640 1 0 $X=373650 $Y=19520
X9361 3 1 137 up_switches<0> BUJI3VX3 $T=379120 24640 1 0 $X=378690 $Y=19520
X9362 3 1 186 7 INJI3VX0 $T=29120 69440 1 0 $X=28690 $Y=64320
X9363 3 1 983 1203 INJI3VX0 $T=39200 69440 1 0 $X=38770 $Y=64320
X9364 3 1 24 200 INJI3VX0 $T=44240 194880 1 180 $X=42130 $Y=194240
X9365 3 1 992 767 INJI3VX0 $T=47040 203840 0 180 $X=44930 $Y=198720
X9366 3 1 979 1422 INJI3VX0 $T=47600 60480 1 0 $X=47170 $Y=55360
X9367 3 1 13 771 INJI3VX0 $T=49840 42560 1 180 $X=47730 $Y=41920
X9368 3 1 10 774 INJI3VX0 $T=49840 42560 0 0 $X=49410 $Y=41920
X9369 3 1 1208 1438 INJI3VX0 $T=52640 60480 1 180 $X=50530 $Y=59840
X9370 3 1 994 998 INJI3VX0 $T=52080 185920 1 0 $X=51650 $Y=180800
X9371 3 1 9 231 INJI3VX0 $T=53200 194880 1 0 $X=52770 $Y=189760
X9372 3 1 244 209 INJI3VX0 $T=57680 33600 1 180 $X=55570 $Y=32960
X9373 3 1 217 202 INJI3VX0 $T=59360 51520 0 180 $X=57250 $Y=46400
X9374 3 1 215 1440 INJI3VX0 $T=59360 96320 1 180 $X=57250 $Y=95680
X9375 3 1 280 205 INJI3VX0 $T=59360 105280 1 180 $X=57250 $Y=104640
X9376 3 1 18 785 INJI3VX0 $T=58240 42560 1 0 $X=57810 $Y=37440
X9377 3 1 218 1414 INJI3VX0 $T=59920 185920 1 0 $X=59490 $Y=180800
X9378 3 1 236 1004 INJI3VX0 $T=63840 176960 1 180 $X=61730 $Y=176320
X9379 3 1 25 1441 INJI3VX0 $T=64400 203840 1 180 $X=62290 $Y=203200
X9380 3 1 1007 1013 INJI3VX0 $T=64400 212800 1 0 $X=63970 $Y=207680
X9381 3 1 232 796 INJI3VX0 $T=68320 203840 1 0 $X=67890 $Y=198720
X9382 3 1 247 1023 INJI3VX0 $T=75040 194880 1 0 $X=74610 $Y=189760
X9383 3 1 283 29 INJI3VX0 $T=81760 105280 0 180 $X=79650 $Y=100160
X9384 3 1 263 1040 INJI3VX0 $T=83440 123200 0 0 $X=83010 $Y=122560
X9385 3 1 274 261 INJI3VX0 $T=85680 194880 1 180 $X=83570 $Y=194240
X9386 3 1 275 805 INJI3VX0 $T=91280 203840 0 180 $X=89170 $Y=198720
X9387 3 1 35 34 INJI3VX0 $T=91840 96320 1 180 $X=89730 $Y=95680
X9388 3 1 281 1220 INJI3VX0 $T=92400 212800 1 0 $X=91970 $Y=207680
X9389 3 1 961 206 INJI3VX0 $T=95200 203840 1 180 $X=93090 $Y=203200
X9390 3 1 823 266 INJI3VX0 $T=96880 176960 1 180 $X=94770 $Y=176320
X9391 3 1 235 286 INJI3VX0 $T=95200 203840 0 0 $X=94770 $Y=203200
X9392 3 1 284 1045 INJI3VX0 $T=98000 105280 1 0 $X=97570 $Y=100160
X9393 3 1 1221 828 INJI3VX0 $T=100240 185920 1 0 $X=99810 $Y=180800
X9394 3 1 826 1397 INJI3VX0 $T=113120 24640 1 0 $X=112690 $Y=19520
X9395 3 1 319 1047 INJI3VX0 $T=124320 194880 0 180 $X=122210 $Y=189760
X9396 3 1 37 1049 INJI3VX0 $T=128800 33600 1 180 $X=126690 $Y=32960
X9397 3 1 833 355 INJI3VX0 $T=133840 194880 0 0 $X=133410 $Y=194240
X9398 3 1 354 838 INJI3VX0 $T=137760 24640 1 180 $X=135650 $Y=24000
X9399 3 1 369 1053 INJI3VX0 $T=137760 194880 1 180 $X=135650 $Y=194240
X9400 3 1 353 843 INJI3VX0 $T=137200 203840 0 0 $X=136770 $Y=203200
X9401 3 1 395 846 INJI3VX0 $T=142800 194880 0 0 $X=142370 $Y=194240
X9402 3 1 385 845 INJI3VX0 $T=149520 33600 1 180 $X=147410 $Y=32960
X9403 3 1 389 849 INJI3VX0 $T=148960 24640 0 0 $X=148530 $Y=24000
X9404 3 1 852 394 INJI3VX0 $T=151760 194880 0 0 $X=151330 $Y=194240
X9405 3 1 368 60 INJI3VX0 $T=155120 203840 1 180 $X=153010 $Y=203200
X9406 3 1 1304 1231 INJI3VX0 $T=155680 185920 1 0 $X=155250 $Y=180800
X9407 3 1 857 1062 INJI3VX0 $T=159600 24640 1 180 $X=157490 $Y=24000
X9408 3 1 856 1064 INJI3VX0 $T=157920 203840 1 0 $X=157490 $Y=198720
X9409 3 1 425 1072 INJI3VX0 $T=163520 24640 0 0 $X=163090 $Y=24000
X9410 3 1 426 420 INJI3VX0 $T=166320 194880 1 180 $X=164210 $Y=194240
X9411 3 1 442 1073 INJI3VX0 $T=171920 194880 1 180 $X=169810 $Y=194240
X9412 3 1 61 867 INJI3VX0 $T=175280 24640 0 0 $X=174850 $Y=24000
X9413 3 1 75 1075 INJI3VX0 $T=182000 194880 1 180 $X=179890 $Y=194240
X9414 3 1 870 1398 INJI3VX0 $T=184240 33600 0 180 $X=182130 $Y=28480
X9415 3 1 464 246 INJI3VX0 $T=184240 194880 0 180 $X=182130 $Y=189760
X9416 3 1 457 1399 INJI3VX0 $T=188160 24640 0 180 $X=186050 $Y=19520
X9417 3 1 1079 448 INJI3VX0 $T=188720 203840 0 180 $X=186610 $Y=198720
X9418 3 1 473 77 INJI3VX0 $T=190960 212800 0 0 $X=190530 $Y=212160
X9419 3 1 474 1237 INJI3VX0 $T=193760 212800 0 0 $X=193330 $Y=212160
X9420 3 1 873 1400 INJI3VX0 $T=198240 33600 1 180 $X=196130 $Y=32960
X9421 3 1 880 1401 INJI3VX0 $T=201040 24640 0 180 $X=198930 $Y=19520
X9422 3 1 94 86 INJI3VX0 $T=201040 203840 0 180 $X=198930 $Y=198720
X9423 3 1 489 882 INJI3VX0 $T=201040 203840 1 0 $X=200610 $Y=198720
X9424 3 1 1084 878 INJI3VX0 $T=204400 203840 0 180 $X=202290 $Y=198720
X9425 3 1 887 1309 INJI3VX0 $T=218960 42560 1 0 $X=218530 $Y=37440
X9426 3 1 101 884 INJI3VX0 $T=221200 24640 1 180 $X=219090 $Y=24000
X9427 3 1 510 1090 INJI3VX0 $T=221200 42560 1 0 $X=220770 $Y=37440
X9428 3 1 507 506 INJI3VX0 $T=227360 185920 1 180 $X=225250 $Y=185280
X9429 3 1 1098 1095 INJI3VX0 $T=233520 24640 1 180 $X=231410 $Y=24000
X9430 3 1 520 103 INJI3VX0 $T=236880 203840 1 180 $X=234770 $Y=203200
X9431 3 1 549 1372 INJI3VX0 $T=240240 194880 0 180 $X=238130 $Y=189760
X9432 3 1 522 895 INJI3VX0 $T=240240 194880 1 0 $X=239810 $Y=189760
X9433 3 1 542 1420 INJI3VX0 $T=246960 194880 1 0 $X=246530 $Y=189760
X9434 3 1 896 1402 INJI3VX0 $T=248640 33600 1 0 $X=248210 $Y=28480
X9435 3 1 897 899 INJI3VX0 $T=250880 42560 0 0 $X=250450 $Y=41920
X9436 3 1 124 1318 INJI3VX0 $T=266000 42560 1 0 $X=265570 $Y=37440
X9437 3 1 595 1255 INJI3VX0 $T=272160 33600 1 0 $X=271730 $Y=28480
X9438 3 1 enable 48 INJI3VX0 $T=276080 185920 0 0 $X=275650 $Y=185280
X9439 3 1 126 618 INJI3VX0 $T=277760 194880 1 0 $X=277330 $Y=189760
X9440 3 1 620 635 INJI3VX0 $T=281120 221760 1 0 $X=280690 $Y=216640
X9441 3 1 910 1403 INJI3VX0 $T=286160 33600 0 180 $X=284050 $Y=28480
X9442 3 1 1121 1260 INJI3VX0 $T=287280 42560 1 0 $X=286850 $Y=37440
X9443 3 1 1124 914 INJI3VX0 $T=299600 33600 0 0 $X=299170 $Y=32960
X9444 3 1 912 658 INJI3VX0 $T=301280 185920 0 0 $X=300850 $Y=185280
X9445 3 1 662 1125 INJI3VX0 $T=301280 194880 1 0 $X=300850 $Y=189760
X9446 3 1 1130 921 INJI3VX0 $T=306320 33600 1 0 $X=305890 $Y=28480
X9447 3 1 665 139 INJI3VX0 $T=313600 185920 1 0 $X=313170 $Y=180800
X9448 3 1 1411 134 INJI3VX0 $T=315840 203840 0 180 $X=313730 $Y=198720
X9449 3 1 672 678 INJI3VX0 $T=324800 194880 0 0 $X=324370 $Y=194240
X9450 3 1 1135 1404 INJI3VX0 $T=328160 42560 0 180 $X=326050 $Y=37440
X9451 3 1 701 688 INJI3VX0 $T=328160 194880 1 180 $X=326050 $Y=194240
X9452 3 1 157 927 INJI3VX0 $T=328720 51520 1 0 $X=328290 $Y=46400
X9453 3 1 687 928 INJI3VX0 $T=330960 203840 1 0 $X=330530 $Y=198720
X9454 3 1 1141 1361 INJI3VX0 $T=334320 203840 0 180 $X=332210 $Y=198720
X9455 3 1 1145 1405 INJI3VX0 $T=335440 33600 0 180 $X=333330 $Y=28480
X9456 3 1 155 1278 INJI3VX0 $T=337680 185920 1 0 $X=337250 $Y=180800
X9457 3 1 935 1146 INJI3VX0 $T=337680 194880 1 0 $X=337250 $Y=189760
X9458 3 1 1277 1147 INJI3VX0 $T=338800 42560 1 0 $X=338370 $Y=37440
X9459 3 1 941 703 INJI3VX0 $T=341040 168000 1 180 $X=338930 $Y=167360
X9460 3 1 938 1406 INJI3VX0 $T=341040 24640 1 0 $X=340610 $Y=19520
X9461 3 1 945 943 INJI3VX0 $T=346640 168000 1 180 $X=344530 $Y=167360
X9462 3 1 730 949 INJI3VX0 $T=350560 42560 1 0 $X=350130 $Y=37440
X9463 3 1 1153 706 INJI3VX0 $T=355040 194880 0 180 $X=352930 $Y=189760
X9464 3 1 951 1330 INJI3VX0 $T=356720 176960 0 0 $X=356290 $Y=176320
X9465 3 1 727 971 INJI3VX0 $T=357840 185920 0 0 $X=357410 $Y=185280
X9466 3 1 1288 1157 INJI3VX0 $T=364560 24640 0 0 $X=364130 $Y=24000
X9467 3 1 164 1407 INJI3VX0 $T=370720 33600 0 180 $X=368610 $Y=28480
X9468 3 1 979 1435 983 NA2JI3VX0 $T=36960 69440 1 0 $X=36530 $Y=64320
X9469 3 1 191 981 764 NA2JI3VX0 $T=42000 60480 1 180 $X=39330 $Y=59840
X9470 3 1 1385 980 765 NA2JI3VX0 $T=43680 203840 0 180 $X=41010 $Y=198720
X9471 3 1 202 991 191 NA2JI3VX0 $T=47040 60480 0 180 $X=44370 $Y=55360
X9472 3 1 193 1436 1160 NA2JI3VX0 $T=49840 42560 0 180 $X=47170 $Y=37440
X9473 3 1 1207 1296 765 NA2JI3VX0 $T=50400 203840 0 180 $X=47730 $Y=198720
X9474 3 1 9 992 995 NA2JI3VX0 $T=53200 194880 1 180 $X=50530 $Y=194240
X9475 3 1 222 772 7 NA2JI3VX0 $T=56560 69440 0 180 $X=53890 $Y=64320
X9476 3 1 16 210 1422 NA2JI3VX0 $T=58800 60480 0 180 $X=56130 $Y=55360
X9477 3 1 261 1297 199 NA2JI3VX0 $T=59360 203840 0 180 $X=56690 $Y=198720
X9478 3 1 1010 784 273 NA2JI3VX0 $T=63840 87360 1 180 $X=61170 $Y=86720
X9479 3 1 1215 788 273 NA2JI3VX0 $T=67760 87360 1 180 $X=65090 $Y=86720
X9480 3 1 793 1216 266 NA2JI3VX0 $T=68880 105280 0 180 $X=66210 $Y=100160
X9481 3 1 253 792 273 NA2JI3VX0 $T=71120 87360 1 180 $X=68450 $Y=86720
X9482 3 1 232 803 247 NA2JI3VX0 $T=71120 203840 0 0 $X=70690 $Y=203200
X9483 3 1 1015 239 231 NA2JI3VX0 $T=73920 194880 0 180 $X=71250 $Y=189760
X9484 3 1 1217 802 273 NA2JI3VX0 $T=75600 87360 1 180 $X=72930 $Y=86720
X9485 3 1 242 1027 1023 NA2JI3VX0 $T=73360 185920 1 0 $X=72930 $Y=180800
X9486 3 1 276 1442 273 NA2JI3VX0 $T=77840 96320 1 0 $X=77410 $Y=91200
X9487 3 1 26 1301 266 NA2JI3VX0 $T=85120 114240 1 0 $X=84690 $Y=109120
X9488 3 1 31 815 266 NA2JI3VX0 $T=89600 123200 1 180 $X=86930 $Y=122560
X9489 3 1 282 1437 1038 NA2JI3VX0 $T=90160 212800 1 0 $X=89730 $Y=207680
X9490 3 1 1219 1443 273 NA2JI3VX0 $T=92960 96320 0 180 $X=90290 $Y=91200
X9491 3 1 49 1439 824 NA2JI3VX0 $T=99680 185920 1 180 $X=97010 $Y=185280
X9492 3 1 269 1337 1038 NA2JI3VX0 $T=98560 203840 0 0 $X=98130 $Y=203200
X9493 3 1 826 1374 107 NA2JI3VX0 $T=99680 24640 1 0 $X=99250 $Y=19520
X9494 3 1 1166 1046 55 NA2JI3VX0 $T=102480 24640 0 0 $X=102050 $Y=24000
X9495 3 1 enable 829 275 NA2JI3VX0 $T=102480 203840 0 0 $X=102050 $Y=203200
X9496 3 1 1166 1222 107 NA2JI3VX0 $T=113680 24640 0 0 $X=113250 $Y=24000
X9497 3 1 319 46 1368 NA2JI3VX0 $T=118160 194880 0 180 $X=115490 $Y=189760
X9498 3 1 1047 312 1368 NA2JI3VX0 $T=121520 194880 0 180 $X=118850 $Y=189760
X9499 3 1 316 1225 107 NA2JI3VX0 $T=123200 24640 0 0 $X=122770 $Y=24000
X9500 3 1 319 460 1224 NA2JI3VX0 $T=123200 203840 1 0 $X=122770 $Y=198720
X9501 3 1 316 1426 55 NA2JI3VX0 $T=127120 24640 0 0 $X=126690 $Y=24000
X9502 3 1 37 1226 107 NA2JI3VX0 $T=128800 33600 1 0 $X=128370 $Y=28480
X9503 3 1 835 837 107 NA2JI3VX0 $T=133280 24640 0 0 $X=132850 $Y=24000
X9504 3 1 348 1052 1444 NA2JI3VX0 $T=134960 203840 1 0 $X=134530 $Y=198720
X9505 3 1 835 1427 55 NA2JI3VX0 $T=135520 33600 1 0 $X=135090 $Y=28480
X9506 3 1 1055 377 355 NA2JI3VX0 $T=136640 185920 1 0 $X=136210 $Y=180800
X9507 3 1 354 841 107 NA2JI3VX0 $T=138320 24640 0 0 $X=137890 $Y=24000
X9508 3 1 350 383 1053 NA2JI3VX0 $T=138320 185920 0 0 $X=137890 $Y=185280
X9509 3 1 839 1054 1444 NA2JI3VX0 $T=138320 203840 1 0 $X=137890 $Y=198720
X9510 3 1 1056 962 107 NA2JI3VX0 $T=139440 33600 0 0 $X=139010 $Y=32960
X9511 3 1 374 1227 107 NA2JI3VX0 $T=141680 24640 0 0 $X=141250 $Y=24000
X9512 3 1 1056 1428 55 NA2JI3VX0 $T=143360 33600 0 0 $X=142930 $Y=32960
X9513 3 1 377 1303 1419 NA2JI3VX0 $T=146160 185920 1 0 $X=145730 $Y=180800
X9514 3 1 385 400 107 NA2JI3VX0 $T=150640 33600 0 0 $X=150210 $Y=32960
X9515 3 1 410 1230 107 NA2JI3VX0 $T=154000 24640 0 0 $X=153570 $Y=24000
X9516 3 1 854 1304 394 NA2JI3VX0 $T=156240 194880 0 180 $X=153570 $Y=189760
X9517 3 1 856 1229 59 NA2JI3VX0 $T=154000 194880 0 0 $X=153570 $Y=194240
X9518 3 1 1068 1233 107 NA2JI3VX0 $T=162960 33600 1 0 $X=162530 $Y=28480
X9519 3 1 419 858 420 NA2JI3VX0 $T=164640 185920 1 0 $X=164210 $Y=180800
X9520 3 1 1070 430 107 NA2JI3VX0 $T=165200 24640 0 0 $X=164770 $Y=24000
X9521 3 1 1073 861 368 NA2JI3VX0 $T=170240 194880 1 180 $X=167570 $Y=194240
X9522 3 1 461 413 1073 NA2JI3VX0 $T=168560 185920 1 0 $X=168130 $Y=180800
X9523 3 1 869 1076 107 NA2JI3VX0 $T=179200 33600 0 0 $X=178770 $Y=32960
X9524 3 1 453 1078 107 NA2JI3VX0 $T=185360 24640 1 180 $X=182690 $Y=24000
X9525 3 1 474 484 473 NA2JI3VX0 $T=187040 212800 0 0 $X=186610 $Y=212160
X9526 3 1 874 1369 107 NA2JI3VX0 $T=197120 42560 0 180 $X=194450 $Y=37440
X9527 3 1 1308 1083 107 NA2JI3VX0 $T=198800 24640 1 180 $X=196130 $Y=24000
X9528 3 1 874 1085 55 NA2JI3VX0 $T=201040 42560 1 0 $X=200610 $Y=37440
X9529 3 1 873 879 107 NA2JI3VX0 $T=201600 33600 0 0 $X=201170 $Y=32960
X9530 3 1 509 477 878 NA2JI3VX0 $T=205520 194880 1 0 $X=205090 $Y=189760
X9531 3 1 511 1312 107 NA2JI3VX0 $T=210560 24640 1 180 $X=207890 $Y=24000
X9532 3 1 1092 1087 107 NA2JI3VX0 $T=210560 33600 1 180 $X=207890 $Y=32960
X9533 3 1 101 1314 107 NA2JI3VX0 $T=221760 33600 1 0 $X=221330 $Y=28480
X9534 3 1 885 1091 508 NA2JI3VX0 $T=225680 203840 1 180 $X=223010 $Y=203200
X9535 3 1 511 1430 490 NA2JI3VX0 $T=225120 24640 0 0 $X=224690 $Y=24000
X9536 3 1 1092 888 490 NA2JI3VX0 $T=225680 33600 0 0 $X=225250 $Y=32960
X9537 3 1 507 1352 885 NA2JI3VX0 $T=227920 203840 1 180 $X=225250 $Y=203200
X9538 3 1 887 1241 107 NA2JI3VX0 $T=226240 42560 1 0 $X=225810 $Y=37440
X9539 3 1 889 1089 107 NA2JI3VX0 $T=232400 42560 0 180 $X=229730 $Y=37440
X9540 3 1 1097 1240 107 NA2JI3VX0 $T=232960 24640 0 180 $X=230290 $Y=19520
X9541 3 1 510 1245 107 NA2JI3VX0 $T=232400 33600 0 0 $X=231970 $Y=32960
X9542 3 1 533 1371 1246 NA2JI3VX0 $T=233520 203840 1 0 $X=233090 $Y=198720
X9543 3 1 889 1099 490 NA2JI3VX0 $T=236320 42560 0 180 $X=233650 $Y=37440
X9544 3 1 1097 1431 490 NA2JI3VX0 $T=234640 24640 1 0 $X=234210 $Y=19520
X9545 3 1 99 97 506 NA2JI3VX0 $T=238560 194880 0 180 $X=235890 $Y=189760
X9546 3 1 1098 1354 107 NA2JI3VX0 $T=238560 24640 0 0 $X=238130 $Y=24000
X9547 3 1 543 1433 490 NA2JI3VX0 $T=240240 42560 1 0 $X=239810 $Y=37440
X9548 3 1 543 1247 107 NA2JI3VX0 $T=241360 33600 0 0 $X=240930 $Y=32960
X9549 3 1 1410 559 1432 NA2JI3VX0 $T=245840 203840 1 0 $X=245410 $Y=198720
X9550 3 1 896 1355 107 NA2JI3VX0 $T=248080 42560 1 0 $X=247650 $Y=37440
X9551 3 1 553 549 1420 NA2JI3VX0 $T=252000 194880 0 180 $X=249330 $Y=189760
X9552 3 1 898 1103 107 NA2JI3VX0 $T=252000 42560 1 0 $X=251570 $Y=37440
X9553 3 1 897 1316 107 NA2JI3VX0 $T=254240 42560 0 0 $X=253810 $Y=41920
X9554 3 1 898 1317 490 NA2JI3VX0 $T=258160 42560 0 180 $X=255490 $Y=37440
X9555 3 1 582 1108 490 NA2JI3VX0 $T=262640 42560 0 180 $X=259970 $Y=37440
X9556 3 1 124 1110 107 NA2JI3VX0 $T=263760 33600 1 180 $X=261090 $Y=32960
X9557 3 1 582 1253 107 NA2JI3VX0 $T=263760 33600 0 0 $X=263330 $Y=32960
X9558 3 1 592 1109 122 NA2JI3VX0 $T=263760 150080 0 0 $X=263330 $Y=149440
X9559 3 1 902 1111 130 NA2JI3VX0 $T=269360 33600 0 0 $X=268930 $Y=32960
X9560 3 1 1118 1117 1115 NA2JI3VX0 $T=280000 203840 0 180 $X=277330 $Y=198720
X9561 3 1 1258 1320 130 NA2JI3VX0 $T=278880 33600 0 0 $X=278450 $Y=32960
X9562 3 1 629 1259 130 NA2JI3VX0 $T=295120 33600 1 180 $X=292450 $Y=32960
X9563 3 1 637 1262 130 NA2JI3VX0 $T=299040 33600 1 180 $X=296370 $Y=32960
X9564 3 1 1127 654 1125 NA2JI3VX0 $T=300720 185920 1 0 $X=300290 $Y=180800
X9565 3 1 915 1265 130 NA2JI3VX0 $T=304080 33600 0 0 $X=303650 $Y=32960
X9566 3 1 662 926 667 NA2JI3VX0 $T=310800 185920 1 0 $X=310370 $Y=180800
X9567 3 1 693 1378 130 NA2JI3VX0 $T=316400 33600 1 180 $X=313730 $Y=32960
X9568 3 1 691 147 130 NA2JI3VX0 $T=325360 51520 1 0 $X=324930 $Y=46400
X9569 3 1 931 682 928 NA2JI3VX0 $T=325360 185920 0 0 $X=324930 $Y=185280
X9570 3 1 142 1324 968 NA2JI3VX0 $T=327600 203840 0 180 $X=324930 $Y=198720
X9571 3 1 687 1271 1272 NA2JI3VX0 $T=328160 194880 0 0 $X=327730 $Y=194240
X9572 3 1 682 930 1137 NA2JI3VX0 $T=329280 185920 1 0 $X=328850 $Y=180800
X9573 3 1 932 969 130 NA2JI3VX0 $T=330400 33600 0 0 $X=329970 $Y=32960
X9574 3 1 158 1379 130 NA2JI3VX0 $T=333760 33600 0 180 $X=331090 $Y=28480
X9575 3 1 160 1326 130 NA2JI3VX0 $T=335440 42560 1 0 $X=335010 $Y=37440
X9576 3 1 701 970 1272 NA2JI3VX0 $T=337680 203840 0 180 $X=335010 $Y=198720
X9577 3 1 713 155 1146 NA2JI3VX0 $T=341040 185920 1 180 $X=338370 $Y=185280
X9578 3 1 944 941 943 NA2JI3VX0 $T=344400 168000 1 180 $X=341730 $Y=167360
X9579 3 1 951 942 1150 NA2JI3VX0 $T=346640 185920 1 180 $X=343970 $Y=185280
X9580 3 1 727 1281 1279 NA2JI3VX0 $T=346080 194880 0 0 $X=345650 $Y=194240
X9581 3 1 165 1282 130 NA2JI3VX0 $T=350000 42560 0 180 $X=347330 $Y=37440
X9582 3 1 167 696 729 NA2JI3VX0 $T=351120 176960 0 180 $X=348450 $Y=171840
X9583 3 1 952 735 130 NA2JI3VX0 $T=357840 24640 0 0 $X=357410 $Y=24000
X9584 3 1 1412 1289 130 NA2JI3VX0 $T=359520 33600 0 0 $X=359090 $Y=32960
X9585 3 1 1155 167 971 NA2JI3VX0 $T=365120 176960 0 180 $X=362450 $Y=171840
X9586 3 1 24 975 195 204 1294 AO22JI3VX1 $T=31360 105280 0 180 $X=25890 $Y=100160
X9587 3 1 973 24 195 179 176 AO22JI3VX1 $T=28560 132160 1 0 $X=28130 $Y=127040
X9588 3 1 972 24 195 5 177 AO22JI3VX1 $T=29120 150080 1 0 $X=28690 $Y=144960
X9589 3 1 761 24 195 1334 178 AO22JI3VX1 $T=29120 168000 0 0 $X=28690 $Y=167360
X9590 3 1 24 760 195 182 763 AO22JI3VX1 $T=29680 114240 0 0 $X=29250 $Y=113600
X9591 3 1 24 183 195 8 181 AO22JI3VX1 $T=33040 105280 1 0 $X=32610 $Y=100160
X9592 3 1 1445 24 195 228 189 AO22JI3VX1 $T=45360 185920 1 180 $X=39890 $Y=185280
X9593 3 1 1446 24 195 9 762 AO22JI3VX1 $T=45360 194880 0 180 $X=39890 $Y=189760
X9594 3 1 1206 24 195 218 188 AO22JI3VX1 $T=47040 176960 0 180 $X=41570 $Y=171840
X9595 3 1 779 235 206 197 187 AO22JI3VX1 $T=49280 159040 0 180 $X=43810 $Y=153920
X9596 3 1 1212 235 206 198 769 AO22JI3VX1 $T=49840 141120 1 180 $X=44370 $Y=140480
X9597 3 1 1295 235 206 773 776 AO22JI3VX1 $T=45920 168000 1 0 $X=45490 $Y=162880
X9598 3 1 235 1159 206 11 988 AO22JI3VX1 $T=52640 123200 1 180 $X=47170 $Y=122560
X9599 3 1 235 15 206 20 989 AO22JI3VX1 $T=55440 123200 0 180 $X=49970 $Y=118080
X9600 3 1 1007 1441 235 1418 207 AO22JI3VX1 $T=61600 203840 1 180 $X=56130 $Y=203200
X9601 3 1 1002 235 206 237 787 AO22JI3VX1 $T=57680 150080 0 0 $X=57250 $Y=149440
X9602 3 1 235 17 206 782 1214 AO22JI3VX1 $T=58240 123200 1 0 $X=57810 $Y=118080
X9603 3 1 235 23 206 793 226 AO22JI3VX1 $T=70560 123200 0 180 $X=65090 $Y=118080
X9604 3 1 1001 24 195 795 243 AO22JI3VX1 $T=69440 141120 0 0 $X=69010 $Y=140480
X9605 3 1 24 249 195 256 238 AO22JI3VX1 $T=78960 114240 0 180 $X=73490 $Y=109120
X9606 3 1 801 235 206 26 291 AO22JI3VX1 $T=73920 123200 0 0 $X=73490 $Y=122560
X9607 3 1 799 235 206 31 285 AO22JI3VX1 $T=74480 150080 1 0 $X=74050 $Y=144960
X9608 3 1 798 24 195 263 255 AO22JI3VX1 $T=76160 141120 0 0 $X=75730 $Y=140480
X9609 3 1 1028 235 206 265 268 AO22JI3VX1 $T=76160 203840 0 0 $X=75730 $Y=203200
X9610 3 1 451 252 805 enable 195 AO22JI3VX1 $T=83440 194880 1 180 $X=77970 $Y=194240
X9611 3 1 1022 24 195 270 290 AO22JI3VX1 $T=79520 114240 1 0 $X=79090 $Y=109120
X9612 3 1 332 368 362 833 320 AO22JI3VX1 $T=128240 203840 1 180 $X=122770 $Y=203200
X9613 3 1 451 1050 314 enable 362 AO22JI3VX1 $T=123760 194880 0 0 $X=123330 $Y=194240
X9614 3 1 410 76 107 857 1065 AO22JI3VX1 $T=156240 33600 1 0 $X=155810 $Y=28480
X9615 3 1 1068 76 107 425 632 AO22JI3VX1 $T=167440 33600 1 0 $X=167010 $Y=28480
X9616 3 1 1070 76 107 61 644 AO22JI3VX1 $T=170240 24640 0 0 $X=169810 $Y=24000
X9617 3 1 869 76 107 870 650 AO22JI3VX1 $T=180880 42560 1 0 $X=180450 $Y=37440
X9618 3 1 453 76 107 457 663 AO22JI3VX1 $T=187600 24640 0 0 $X=187170 $Y=24000
X9619 3 1 1308 649 107 880 478 AO22JI3VX1 $T=201600 24640 0 0 $X=201170 $Y=24000
X9620 3 1 483 86 882 474 475 AO22JI3VX1 $T=208880 203840 1 180 $X=203410 $Y=203200
X9621 3 1 1088 86 882 1084 883 AO22JI3VX1 $T=204960 203840 1 0 $X=204530 $Y=198720
X9622 3 1 507 508 86 1350 886 AO22JI3VX1 $T=225120 203840 0 180 $X=219650 $Y=198720
X9623 3 1 902 649 130 595 680 AO22JI3VX1 $T=272160 33600 0 0 $X=271730 $Y=32960
X9624 3 1 637 649 130 1124 137 AO22JI3VX1 $T=297920 42560 1 0 $X=297490 $Y=37440
X9625 3 1 915 649 130 1130 704 AO22JI3VX1 $T=308000 33600 0 0 $X=307570 $Y=32960
X9626 3 1 925 672 968 665 144 AO22JI3VX1 $T=316960 194880 0 180 $X=311490 $Y=189760
X9627 3 1 693 649 130 1135 150 AO22JI3VX1 $T=324800 33600 0 0 $X=324370 $Y=32960
X9628 3 1 691 649 130 157 1139 AO22JI3VX1 $T=325920 42560 0 0 $X=325490 $Y=41920
X9629 3 1 932 649 130 1145 736 AO22JI3VX1 $T=335440 33600 1 0 $X=335010 $Y=28480
X9630 3 1 672 934 935 48 715 AO22JI3VX1 $T=336000 194880 0 0 $X=335570 $Y=194240
X9631 3 1 158 649 130 938 719 AO22JI3VX1 $T=341600 33600 1 0 $X=341170 $Y=28480
X9632 3 1 160 649 130 1277 946 AO22JI3VX1 $T=341600 42560 1 0 $X=341170 $Y=37440
X9633 3 1 672 1373 1279 1283 1197 AO22JI3VX1 $T=348880 194880 0 0 $X=348450 $Y=194240
X9634 3 1 1447 672 945 48 743 AO22JI3VX1 $T=350560 176960 0 0 $X=350130 $Y=176320
X9635 3 1 1151 672 951 48 1290 AO22JI3VX1 $T=350560 185920 0 0 $X=350130 $Y=185280
X9636 3 1 1412 649 130 164 1152 AO22JI3VX1 $T=357840 33600 1 180 $X=352370 $Y=32960
X9637 3 1 952 649 130 1288 1284 AO22JI3VX1 $T=358400 33600 0 180 $X=352930 $Y=28480
X9638 3 1 165 649 130 730 947 AO22JI3VX1 $T=358400 42560 0 180 $X=352930 $Y=37440
X9639 3 1 673 1269 668 660 1187 OR4JI3VX2 $T=316960 24640 1 180 $X=309250 $Y=24000
X9640 3 1 434 56 INJI3VX2 $T=173600 168000 1 0 $X=173170 $Y=162880
X9641 3 1 434 71 INJI3VX2 $T=177520 185920 0 0 $X=177090 $Y=185280
X9642 3 1 113 600 INJI3VX2 $T=223440 221760 1 0 $X=223010 $Y=216640
X9643 3 1 107 768 196 1202 AO21JI3VX1 $T=43120 78400 1 180 $X=38210 $Y=77760
X9644 3 1 24 992 195 765 AO21JI3VX1 $T=49840 194880 1 180 $X=44930 $Y=194240
X9645 3 1 247 206 800 1011 AO21JI3VX1 $T=73360 212800 0 180 $X=68450 $Y=207680
X9646 3 1 818 1040 284 1302 AO21JI3VX1 $T=92400 114240 0 180 $X=87490 $Y=109120
X9647 3 1 843 368 362 1444 AO21JI3VX1 $T=145040 203840 0 180 $X=140130 $Y=198720
X9648 3 1 48 642 1123 1122 AO21JI3VX1 $T=296800 194880 0 180 $X=291890 $Y=189760
X9649 3 1 227 1009 278 NO2I1JI3VX1 $T=64960 194880 0 0 $X=64530 $Y=194240
X9650 3 1 1027 250 1415 NO2I1JI3VX1 $T=77840 176960 1 180 $X=74050 $Y=176320
X9651 3 1 323 1019 256 NO2I1JI3VX1 $T=80080 96320 1 180 $X=76290 $Y=95680
X9652 3 1 33 296 270 NO2I1JI3VX1 $T=86800 105280 0 0 $X=86370 $Y=104640
X9653 3 1 272 817 282 NO2I1JI3VX1 $T=88480 185920 0 0 $X=88050 $Y=185280
X9654 3 1 278 821 1041 NO2I1JI3VX1 $T=91840 194880 0 0 $X=91410 $Y=194240
X9655 3 1 1224 275 319 NO2I1JI3VX1 $T=122080 203840 0 180 $X=118290 $Y=198720
X9656 3 1 308 1224 38 NO2I1JI3VX1 $T=123200 194880 1 180 $X=119410 $Y=194240
X9657 3 1 348 54 834 NO2I1JI3VX1 $T=128800 185920 0 0 $X=128370 $Y=185280
X9658 3 1 346 351 54 NO2I1JI3VX1 $T=134400 194880 1 0 $X=133970 $Y=189760
X9659 3 1 861 868 362 NO2I1JI3VX1 $T=166880 203840 1 0 $X=166450 $Y=198720
X9660 3 1 79 1417 474 NO2I1JI3VX1 $T=196560 194880 0 0 $X=196130 $Y=194240
X9661 3 1 98 482 885 NO2I1JI3VX1 $T=222320 185920 1 180 $X=218530 $Y=185280
X9662 3 1 122 1113 592 NO2I1JI3VX1 $T=267120 150080 0 0 $X=266690 $Y=149440
X9663 3 1 654 917 1131 NO2I1JI3VX1 $T=306320 176960 1 180 $X=302530 $Y=176320
X9664 3 1 235 959 796 247 NA3JI3VX0 $T=70000 194880 0 0 $X=69570 $Y=194240
X9665 3 1 802 1014 1396 1216 NA3JI3VX0 $T=74480 96320 1 180 $X=71250 $Y=95680
X9666 3 1 259 808 807 272 NA3JI3VX0 $T=81200 185920 1 0 $X=80770 $Y=180800
X9667 3 1 1442 1030 809 1301 NA3JI3VX0 $T=83440 96320 1 0 $X=83010 $Y=91200
X9668 3 1 279 36 277 272 NA3JI3VX0 $T=85680 185920 1 0 $X=85250 $Y=180800
X9669 3 1 1443 1036 816 815 NA3JI3VX0 $T=89600 96320 0 180 $X=86370 $Y=91200
X9670 3 1 1047 314 308 38 NA3JI3VX0 $T=115920 194880 0 0 $X=115490 $Y=194240
X9671 3 1 424 405 383 1168 NA3JI3VX0 $T=149520 194880 0 180 $X=146290 $Y=189760
X9672 3 1 1061 313 1448 1059 NA3JI3VX0 $T=155120 185920 1 180 $X=151890 $Y=185280
X9673 3 1 351 1376 413 417 NA3JI3VX0 $T=160160 194880 1 0 $X=159730 $Y=189760
X9674 3 1 859 409 1448 858 NA3JI3VX0 $T=164080 185920 1 180 $X=160850 $Y=185280
X9675 3 1 1449 1173 858 860 NA3JI3VX0 $T=167440 185920 1 180 $X=164210 $Y=185280
X9676 3 1 1429 859 860 417 NA3JI3VX0 $T=167440 194880 0 180 $X=164210 $Y=189760
X9677 3 1 368 1234 448 442 NA3JI3VX0 $T=172480 194880 0 0 $X=172050 $Y=194240
X9678 3 1 1079 63 442 75 NA3JI3VX0 $T=179200 194880 1 180 $X=175970 $Y=194240
X9679 3 1 1377 156 923 132 NA3JI3VX0 $T=310800 176960 1 0 $X=310370 $Y=171840
X9680 3 1 672 1266 134 642 NA3JI3VX0 $T=313600 194880 1 180 $X=310370 $Y=194240
X9681 3 1 676 924 697 923 NA3JI3VX0 $T=316960 176960 0 180 $X=313730 $Y=171840
X9682 3 1 156 1325 1134 697 NA3JI3VX0 $T=333200 176960 0 0 $X=332770 $Y=176320
X9683 3 1 107 196 982 OR2JI3VX0 $T=43120 69440 1 180 $X=39330 $Y=68800
X9684 3 1 191 202 957 OR2JI3VX0 $T=41440 60480 1 0 $X=41010 $Y=55360
X9685 3 1 1013 794 1020 OR2JI3VX0 $T=69440 185920 0 0 $X=69010 $Y=185280
X9686 3 1 803 1013 1031 OR2JI3VX0 $T=74480 203840 1 0 $X=74050 $Y=198720
X9687 3 1 1053 350 1168 OR2JI3VX0 $T=138320 194880 1 0 $X=137890 $Y=189760
X9688 3 1 420 419 860 OR2JI3VX0 $T=161280 185920 1 0 $X=160850 $Y=180800
X9689 3 1 1075 439 417 OR2JI3VX0 $T=180880 194880 0 180 $X=177090 $Y=189760
X9690 3 1 460 48 447 OR2JI3VX0 $T=184800 185920 1 180 $X=181010 $Y=185280
X9691 3 1 1237 872 876 OR2JI3VX0 $T=193200 194880 0 0 $X=192770 $Y=194240
X9692 3 1 103 1101 1353 OR2JI3VX0 $T=235760 185920 0 180 $X=231970 $Y=180800
X9693 3 1 1125 1127 132 OR2JI3VX0 $T=296800 176960 0 0 $X=296370 $Y=176320
X9694 3 1 940 706 937 OR2JI3VX0 $T=343280 194880 0 180 $X=339490 $Y=189760
X9695 3 1 enable 1341 49 260 1223 AO211JI3VX1 $T=113120 185920 0 0 $X=112690 $Y=185280
X9696 3 1 761 234 184 978 HAJI3VX1 $T=28000 159040 0 0 $X=27570 $Y=158400
X9697 3 1 1295 234 201 987 HAJI3VX1 $T=48160 159040 1 180 $X=39890 $Y=158400
X9698 3 1 1206 208 218 994 HAJI3VX1 $T=44800 176960 0 0 $X=44370 $Y=176320
X9699 3 1 1445 228 994 995 HAJI3VX1 $T=45920 185920 0 0 $X=45490 $Y=185280
X9700 3 1 332 833 836 353 HAJI3VX1 $T=126000 203840 1 0 $X=125570 $Y=198720
X9701 3 1 1119 624 1450 1115 HAJI3VX1 $T=281120 203840 1 0 $X=280690 $Y=198720
X9702 3 1 634 630 1321 1450 HAJI3VX1 $T=296800 203840 0 180 $X=288530 $Y=198720
X9703 3 1 1447 945 1149 1150 HAJI3VX1 $T=349440 176960 1 180 $X=341170 $Y=176320
X9704 3 1 813 820 821 292 OA21JI3VX1 $T=91280 194880 1 0 $X=90850 $Y=189760
X9705 3 1 1117 1115 906 1112 OA21JI3VX1 $T=276640 203840 0 180 $X=271730 $Y=198720
X9706 3 1 9 995 1446 EO2JI3VX0 $T=52080 194880 0 180 $X=46050 $Y=189760
X9707 3 1 1024 283 1035 EO2JI3VX0 $T=81760 105280 1 0 $X=81330 $Y=100160
X9708 3 1 284 825 960 EO2JI3VX0 $T=96880 105280 0 180 $X=90850 $Y=100160
X9709 3 1 583 IC_addr<1> 1106 EO2JI3VX0 $T=250880 212800 0 0 $X=250450 $Y=212160
X9710 3 1 1104 IC_addr<0> 901 EO2JI3VX0 $T=253120 221760 1 0 $X=252690 $Y=216640
X9711 3 1 951 1150 1151 EO2JI3VX0 $T=345520 185920 1 0 $X=345090 $Y=180800
X9712 3 1 808 824 812 1218 NO3JI3VX0 $T=84560 185920 0 0 $X=84130 $Y=185280
X9713 3 1 1416 273 1221 260 NO3JI3VX0 $T=101360 176960 1 180 $X=97570 $Y=176320
X9714 3 1 387 1059 1419 851 NO3JI3VX0 $T=148400 185920 1 0 $X=147970 $Y=180800
X9715 3 1 405 1061 1376 1173 NO3JI3VX0 $T=156800 194880 1 0 $X=156370 $Y=189760
X9716 3 1 1236 1082 482 79 NO3JI3VX0 $T=196000 185920 1 180 $X=192210 $Y=185280
X9717 3 1 1106 122 901 593 NO3JI3VX0 $T=259840 203840 0 0 $X=259410 $Y=203200
X9718 3 1 1137 1360 1144 690 NO3JI3VX0 $T=330960 185920 1 180 $X=327170 $Y=185280
X9719 3 1 939 936 162 48 NO3JI3VX0 $T=342160 176960 0 180 $X=338370 $Y=171840
X9720 3 1 817 277 279 819 274 AN31JI3VX1 $T=90720 185920 1 0 $X=90290 $Y=180800
X9721 3 1 1384 1082 515 260 447 AN31JI3VX1 $T=189840 185920 1 180 $X=185490 $Y=185280
X9722 3 1 1413 991 768 AND2JI3VX0 $T=48160 69440 0 180 $X=44370 $Y=64320
X9723 3 1 388 395 836 AND2JI3VX0 $T=142800 194880 1 180 $X=139010 $Y=194240
X9724 3 1 77 872 79 AND2JI3VX0 $T=193200 194880 0 180 $X=189410 $Y=189760
X9725 3 1 103 1101 516 AND2JI3VX0 $T=239120 185920 0 180 $X=235330 $Y=180800
X9726 3 1 620 617 1321 AND2JI3VX0 $T=291760 212800 0 180 $X=287970 $Y=207680
X9727 3 1 1244 515 892 1394 NO3I1JI3VX1 $T=236880 185920 1 180 $X=231970 $Y=185280
X9728 3 1 1063 1064 1448 1231 403 AN211JI3VX1 $T=160160 185920 1 180 $X=155250 $Y=185280
X9729 3 1 1274 139 1134 703 718 AN211JI3VX1 $T=335440 168000 1 180 $X=330530 $Y=167360
X9730 3 1 714 706 1136 1278 153 AN211JI3VX1 $T=340480 176960 1 180 $X=335570 $Y=176320
X9731 3 1 1073 461 1449 866 NO22JI3VX1 $T=168560 185920 0 0 $X=168130 $Y=185280
X9732 3 1 577 43 1113 NA2JI3VX2 $T=275520 150080 0 180 $X=271170 $Y=144960
X9733 3 1 577 1109 307 NO2JI3VX2 $T=259280 150080 0 0 $X=258850 $Y=149440
X9734 3 1 1109 44 577 NA2I1JI3VX2 $T=262080 150080 1 0 $X=261650 $Y=144960
X9735 3 1 577 45 1113 NA2I1JI3VX2 $T=273280 150080 0 0 $X=272850 $Y=149440
X9736 3 1 DECAP25JI3V $T=20160 24640 1 0 $X=19730 $Y=19520
X9737 3 1 DECAP25JI3V $T=20160 24640 0 0 $X=19730 $Y=24000
X9738 3 1 DECAP25JI3V $T=20160 87360 0 0 $X=19730 $Y=86720
X9739 3 1 DECAP25JI3V $T=20160 168000 1 0 $X=19730 $Y=162880
X9740 3 1 DECAP25JI3V $T=20160 212800 0 0 $X=19730 $Y=212160
X9741 3 1 DECAP25JI3V $T=20160 221760 1 0 $X=19730 $Y=216640
X9742 3 1 DECAP25JI3V $T=33040 33600 1 0 $X=32610 $Y=28480
X9743 3 1 DECAP25JI3V $T=34160 24640 1 0 $X=33730 $Y=19520
X9744 3 1 DECAP25JI3V $T=34160 87360 0 0 $X=33730 $Y=86720
X9745 3 1 DECAP25JI3V $T=34160 221760 1 0 $X=33730 $Y=216640
X9746 3 1 DECAP25JI3V $T=47040 33600 1 0 $X=46610 $Y=28480
X9747 3 1 DECAP25JI3V $T=99120 123200 0 0 $X=98690 $Y=122560
X9748 3 1 DECAP25JI3V $T=191520 96320 0 0 $X=191090 $Y=95680
X9749 3 1 DECAP25JI3V $T=212240 105280 1 0 $X=211810 $Y=100160
X9750 3 1 DECAP25JI3V $T=213920 114240 1 0 $X=213490 $Y=109120
X9751 3 1 DECAP25JI3V $T=260400 114240 0 0 $X=259970 $Y=113600
X9752 3 1 DECAP25JI3V $T=301280 69440 0 0 $X=300850 $Y=68800
X9753 3 1 DECAP25JI3V $T=309120 132160 0 0 $X=308690 $Y=131520
X9754 3 1 DECAP25JI3V $T=310800 78400 0 0 $X=310370 $Y=77760
X9755 3 1 DECAP25JI3V $T=341040 221760 1 0 $X=340610 $Y=216640
X9756 3 1 DECAP25JI3V $T=344400 212800 0 0 $X=343970 $Y=212160
X9757 3 1 DECAP25JI3V $T=344960 87360 1 0 $X=344530 $Y=82240
X9758 3 1 DECAP25JI3V $T=344960 212800 1 0 $X=344530 $Y=207680
X9759 3 1 DECAP25JI3V $T=355040 221760 1 0 $X=354610 $Y=216640
X9760 3 1 DECAP25JI3V $T=358400 105280 0 0 $X=357970 $Y=104640
X9761 3 1 DECAP25JI3V $T=358400 212800 0 0 $X=357970 $Y=212160
X9762 3 1 DECAP25JI3V $T=358960 87360 1 0 $X=358530 $Y=82240
X9763 3 1 DECAP25JI3V $T=358960 212800 1 0 $X=358530 $Y=207680
X9764 3 1 DECAP25JI3V $T=361760 150080 1 0 $X=361330 $Y=144960
X9765 3 1 DECAP25JI3V $T=362880 203840 0 0 $X=362450 $Y=203200
X9766 3 1 DECAP25JI3V $T=364000 176960 0 0 $X=363570 $Y=176320
X9767 3 1 DECAP25JI3V $T=365120 132160 1 0 $X=364690 $Y=127040
X9768 3 1 DECAP25JI3V $T=366240 24640 0 0 $X=365810 $Y=24000
X9769 3 1 DECAP25JI3V $T=367360 203840 1 0 $X=366930 $Y=198720
X9770 3 1 DECAP25JI3V $T=369040 221760 1 0 $X=368610 $Y=216640
X9771 3 1 DECAP25JI3V $T=371280 194880 0 0 $X=370850 $Y=194240
X9772 3 1 DECAP25JI3V $T=372400 105280 0 0 $X=371970 $Y=104640
X9773 3 1 DECAP25JI3V $T=372400 194880 1 0 $X=371970 $Y=189760
X9774 3 1 DECAP25JI3V $T=372400 212800 0 0 $X=371970 $Y=212160
X9775 3 1 DECAP25JI3V $T=372960 87360 1 0 $X=372530 $Y=82240
X9776 3 1 DECAP25JI3V $T=372960 212800 1 0 $X=372530 $Y=207680
X9777 3 1 DECAP25JI3V $T=374080 185920 1 0 $X=373650 $Y=180800
X9778 3 1 DECAP25JI3V $T=374640 185920 0 0 $X=374210 $Y=185280
X9779 3 1 DECAP25JI3V $T=375200 123200 0 0 $X=374770 $Y=122560
X9780 3 1 DECAP25JI3V $T=375760 150080 1 0 $X=375330 $Y=144960
X9781 3 1 DECAP25JI3V $T=376880 203840 0 0 $X=376450 $Y=203200
X9782 3 1 DECAP25JI3V $T=378000 176960 0 0 $X=377570 $Y=176320
X9783 3 1 DECAP25JI3V $T=378560 78400 0 0 $X=378130 $Y=77760
X9784 3 1 DECAP25JI3V $T=392560 87360 1 180 $X=378130 $Y=86720
X9785 3 1 DECAP25JI3V $T=378560 96320 1 0 $X=378130 $Y=91200
X9786 3 1 DECAP25JI3V $T=378560 150080 0 0 $X=378130 $Y=149440
X9787 3 1 DECAP25JI3V $T=379120 51520 1 0 $X=378690 $Y=46400
X9788 3 1 DECAP25JI3V $T=379120 51520 0 0 $X=378690 $Y=50880
X9789 3 1 DECAP25JI3V $T=379120 60480 1 0 $X=378690 $Y=55360
X9790 3 1 DECAP25JI3V $T=379120 60480 0 0 $X=378690 $Y=59840
X9791 3 1 DECAP25JI3V $T=379120 69440 0 0 $X=378690 $Y=68800
X9792 3 1 DECAP25JI3V $T=379120 132160 1 0 $X=378690 $Y=127040
X9793 3 1 DECAP25JI3V $T=379120 159040 0 0 $X=378690 $Y=158400
X9794 3 1 DECAP25JI3V $T=379120 168000 0 0 $X=378690 $Y=167360
X9795 3 1 DECAP25JI3V $T=379680 33600 0 0 $X=379250 $Y=32960
X9796 3 1 DECAP25JI3V $T=380240 24640 0 0 $X=379810 $Y=24000
X9797 3 1 DECAP25JI3V $T=380240 159040 1 0 $X=379810 $Y=153920
X9798 3 1 DECAP25JI3V $T=380800 33600 1 0 $X=380370 $Y=28480
X9799 3 1 DECAP25JI3V $T=380800 114240 1 0 $X=380370 $Y=109120
X9800 3 1 DECAP25JI3V $T=380800 141120 0 0 $X=380370 $Y=140480
X9801 3 1 DECAP25JI3V $T=381360 203840 1 0 $X=380930 $Y=198720
X9802 3 1 DECAP25JI3V $T=381920 96320 0 0 $X=381490 $Y=95680
X9803 3 1 DECAP25JI3V $T=381920 105280 1 0 $X=381490 $Y=100160
X9804 3 1 DECAP25JI3V $T=381920 114240 0 0 $X=381490 $Y=113600
X9805 3 1 DECAP25JI3V $T=381920 132160 0 0 $X=381490 $Y=131520
X9806 3 1 DECAP25JI3V $T=381920 141120 1 0 $X=381490 $Y=136000
X9807 3 1 DECAP25JI3V $T=382480 69440 1 0 $X=382050 $Y=64320
X9808 3 1 DECAP25JI3V $T=383040 24640 1 0 $X=382610 $Y=19520
X9809 3 1 DECAP25JI3V $T=383040 221760 1 0 $X=382610 $Y=216640
X9810 3 1 DECAP25JI3V $T=385280 194880 0 0 $X=384850 $Y=194240
X9811 3 1 DECAP25JI3V $T=386400 105280 0 0 $X=385970 $Y=104640
X9812 3 1 DECAP25JI3V $T=386400 123200 1 0 $X=385970 $Y=118080
X9813 3 1 DECAP25JI3V $T=386400 194880 1 0 $X=385970 $Y=189760
X9814 3 1 DECAP25JI3V $T=386400 212800 0 0 $X=385970 $Y=212160
X9815 3 1 DECAP25JI3V $T=386960 78400 1 0 $X=386530 $Y=73280
X9816 3 1 DECAP25JI3V $T=386960 87360 1 0 $X=386530 $Y=82240
X9817 3 1 DECAP25JI3V $T=386960 212800 1 0 $X=386530 $Y=207680
X9818 3 1 DECAP25JI3V $T=387520 176960 1 0 $X=387090 $Y=171840
X9819 3 1 DECAP25JI3V $T=388080 185920 1 0 $X=387650 $Y=180800
X9820 3 1 DECAP25JI3V $T=388640 185920 0 0 $X=388210 $Y=185280
X9821 3 1 DECAP25JI3V $T=389200 123200 0 0 $X=388770 $Y=122560
X9822 3 1 DECAP25JI3V $T=389760 150080 1 0 $X=389330 $Y=144960
X9823 3 1 DECAP25JI3V $T=390880 203840 0 0 $X=390450 $Y=203200
X9824 3 1 DECAP25JI3V $T=392000 176960 0 0 $X=391570 $Y=176320
X9825 3 1 DECAP25JI3V $T=392560 78400 0 0 $X=392130 $Y=77760
X9826 3 1 DECAP25JI3V $T=392560 87360 0 0 $X=392130 $Y=86720
X9827 3 1 DECAP25JI3V $T=392560 96320 1 0 $X=392130 $Y=91200
X9828 3 1 DECAP25JI3V $T=392560 150080 0 0 $X=392130 $Y=149440
X9829 3 1 DECAP25JI3V $T=393120 42560 1 0 $X=392690 $Y=37440
X9830 3 1 DECAP25JI3V $T=393120 42560 0 0 $X=392690 $Y=41920
X9831 3 1 DECAP25JI3V $T=393120 51520 1 0 $X=392690 $Y=46400
X9832 3 1 DECAP25JI3V $T=393120 51520 0 0 $X=392690 $Y=50880
X9833 3 1 DECAP25JI3V $T=393120 60480 1 0 $X=392690 $Y=55360
X9834 3 1 DECAP25JI3V $T=393120 60480 0 0 $X=392690 $Y=59840
X9835 3 1 DECAP25JI3V $T=393120 69440 0 0 $X=392690 $Y=68800
X9836 3 1 DECAP25JI3V $T=393120 132160 1 0 $X=392690 $Y=127040
X9837 3 1 DECAP25JI3V $T=393120 159040 0 0 $X=392690 $Y=158400
X9838 3 1 DECAP25JI3V $T=393120 168000 1 0 $X=392690 $Y=162880
X9839 3 1 DECAP25JI3V $T=393120 168000 0 0 $X=392690 $Y=167360
X9840 3 1 DECAP25JI3V $T=393680 33600 0 0 $X=393250 $Y=32960
X9841 3 1 DECAP25JI3V $T=394240 24640 0 0 $X=393810 $Y=24000
X9842 3 1 DECAP25JI3V $T=394240 159040 1 0 $X=393810 $Y=153920
X9843 3 1 DECAP25JI3V $T=394800 33600 1 0 $X=394370 $Y=28480
X9844 3 1 DECAP25JI3V $T=394800 114240 1 0 $X=394370 $Y=109120
X9845 3 1 DECAP25JI3V $T=394800 141120 0 0 $X=394370 $Y=140480
X9846 3 1 DECAP25JI3V $T=395360 203840 1 0 $X=394930 $Y=198720
X9847 3 1 DECAP25JI3V $T=395920 96320 0 0 $X=395490 $Y=95680
X9848 3 1 DECAP25JI3V $T=395920 105280 1 0 $X=395490 $Y=100160
X9849 3 1 DECAP25JI3V $T=395920 114240 0 0 $X=395490 $Y=113600
X9850 3 1 DECAP25JI3V $T=395920 132160 0 0 $X=395490 $Y=131520
X9851 3 1 DECAP25JI3V $T=395920 141120 1 0 $X=395490 $Y=136000
X9852 3 1 DECAP25JI3V $T=396480 69440 1 0 $X=396050 $Y=64320
X9853 3 1 DECAP25JI3V $T=397040 24640 1 0 $X=396610 $Y=19520
X9854 3 1 DECAP25JI3V $T=397040 221760 1 0 $X=396610 $Y=216640
X9855 3 1 DECAP25JI3V $T=399280 194880 0 0 $X=398850 $Y=194240
X9856 3 1 DECAP25JI3V $T=400400 105280 0 0 $X=399970 $Y=104640
X9857 3 1 DECAP25JI3V $T=400400 123200 1 0 $X=399970 $Y=118080
X9858 3 1 DECAP25JI3V $T=400400 194880 1 0 $X=399970 $Y=189760
X9859 3 1 DECAP25JI3V $T=400400 212800 0 0 $X=399970 $Y=212160
X9860 3 1 DECAP25JI3V $T=401520 176960 1 0 $X=401090 $Y=171840
X9861 3 1 DECAP25JI3V $T=402640 185920 0 0 $X=402210 $Y=185280
X9862 3 1 DECAP25JI3V $T=403200 123200 0 0 $X=402770 $Y=122560
X9863 3 1 DECAP25JI3V $T=407120 42560 1 0 $X=406690 $Y=37440
X9864 3 1 DECAP25JI3V $T=407120 42560 0 0 $X=406690 $Y=41920
X9865 3 1 DECAP25JI3V $T=407120 51520 1 0 $X=406690 $Y=46400
X9866 3 1 DECAP25JI3V $T=407120 51520 0 0 $X=406690 $Y=50880
X9867 3 1 DECAP25JI3V $T=407120 60480 1 0 $X=406690 $Y=55360
X9868 3 1 DECAP25JI3V $T=407120 60480 0 0 $X=406690 $Y=59840
X9869 3 1 DECAP25JI3V $T=407120 69440 0 0 $X=406690 $Y=68800
X9870 3 1 DECAP25JI3V $T=407120 132160 1 0 $X=406690 $Y=127040
X9871 3 1 DECAP25JI3V $T=407120 159040 0 0 $X=406690 $Y=158400
X9872 3 1 DECAP25JI3V $T=407120 168000 1 0 $X=406690 $Y=162880
X9873 3 1 DECAP25JI3V $T=407120 168000 0 0 $X=406690 $Y=167360
X9874 3 1 DECAP25JI3V $T=408240 24640 0 0 $X=407810 $Y=24000
X9875 3 1 DECAP25JI3V $T=408240 159040 1 0 $X=407810 $Y=153920
X9876 3 1 DECAP25JI3V $T=411040 24640 1 0 $X=410610 $Y=19520
X9877 3 1 DECAP25JI3V $T=411040 221760 1 0 $X=410610 $Y=216640
X9878 3 1 DECAP10JI3V $T=20160 60480 0 0 $X=19730 $Y=59840
X9879 3 1 DECAP10JI3V $T=20160 69440 1 0 $X=19730 $Y=64320
X9880 3 1 DECAP10JI3V $T=20160 87360 1 0 $X=19730 $Y=82240
X9881 3 1 DECAP10JI3V $T=20160 96320 1 0 $X=19730 $Y=91200
X9882 3 1 DECAP10JI3V $T=20160 168000 0 0 $X=19730 $Y=167360
X9883 3 1 DECAP10JI3V $T=20160 212800 1 0 $X=19730 $Y=207680
X9884 3 1 DECAP10JI3V $T=24080 114240 0 0 $X=23650 $Y=113600
X9885 3 1 DECAP10JI3V $T=39200 141120 0 0 $X=38770 $Y=140480
X9886 3 1 DECAP10JI3V $T=48160 24640 1 0 $X=47730 $Y=19520
X9887 3 1 DECAP10JI3V $T=48160 87360 0 0 $X=47730 $Y=86720
X9888 3 1 DECAP10JI3V $T=48160 221760 1 0 $X=47730 $Y=216640
X9889 3 1 DECAP10JI3V $T=69440 78400 0 180 $X=63410 $Y=73280
X9890 3 1 DECAP10JI3V $T=68320 159040 0 0 $X=67890 $Y=158400
X9891 3 1 DECAP10JI3V $T=100800 176960 1 0 $X=100370 $Y=171840
X9892 3 1 DECAP10JI3V $T=104720 24640 0 0 $X=104290 $Y=24000
X9893 3 1 DECAP10JI3V $T=133280 176960 1 0 $X=132850 $Y=171840
X9894 3 1 DECAP10JI3V $T=148400 96320 1 0 $X=147970 $Y=91200
X9895 3 1 DECAP10JI3V $T=148400 141120 1 0 $X=147970 $Y=136000
X9896 3 1 DECAP10JI3V $T=197680 123200 0 0 $X=197250 $Y=122560
X9897 3 1 DECAP10JI3V $T=197680 132160 0 0 $X=197250 $Y=131520
X9898 3 1 DECAP10JI3V $T=205520 96320 0 0 $X=205090 $Y=95680
X9899 3 1 DECAP10JI3V $T=210000 123200 1 0 $X=209570 $Y=118080
X9900 3 1 DECAP10JI3V $T=210000 159040 1 0 $X=209570 $Y=153920
X9901 3 1 DECAP10JI3V $T=212800 24640 1 0 $X=212370 $Y=19520
X9902 3 1 DECAP10JI3V $T=213360 33600 1 0 $X=212930 $Y=28480
X9903 3 1 DECAP10JI3V $T=226240 105280 1 0 $X=225810 $Y=100160
X9904 3 1 DECAP10JI3V $T=239120 159040 0 0 $X=238690 $Y=158400
X9905 3 1 DECAP10JI3V $T=240240 96320 0 0 $X=239810 $Y=95680
X9906 3 1 DECAP10JI3V $T=246960 141120 1 0 $X=246530 $Y=136000
X9907 3 1 DECAP10JI3V $T=310240 141120 1 0 $X=309810 $Y=136000
X9908 3 1 DECAP10JI3V $T=315280 69440 0 0 $X=314850 $Y=68800
X9909 3 1 DECAP10JI3V $T=315280 87360 1 0 $X=314850 $Y=82240
X9910 3 1 DECAP10JI3V $T=316400 24640 1 0 $X=315970 $Y=19520
X9911 3 1 DECAP10JI3V $T=317520 159040 1 0 $X=317090 $Y=153920
X9912 3 1 DECAP10JI3V $T=317520 194880 0 0 $X=317090 $Y=194240
X9913 3 1 DECAP10JI3V $T=317520 203840 0 0 $X=317090 $Y=203200
X9914 3 1 DECAP10JI3V $T=318080 24640 0 0 $X=317650 $Y=24000
X9915 3 1 DECAP10JI3V $T=338800 159040 0 0 $X=338370 $Y=158400
X9916 3 1 DECAP10JI3V $T=351680 105280 1 0 $X=351250 $Y=100160
X9917 3 1 DECAP10JI3V $T=353360 96320 0 0 $X=352930 $Y=95680
X9918 3 1 DECAP10JI3V $T=403760 150080 1 0 $X=403330 $Y=144960
X9919 3 1 DECAP10JI3V $T=407680 33600 0 0 $X=407250 $Y=32960
X9920 3 1 DECAP10JI3V $T=415520 176960 1 0 $X=415090 $Y=171840
X9921 3 1 DECAP7JI3V $T=20160 33600 0 0 $X=19730 $Y=32960
X9922 3 1 DECAP7JI3V $T=20160 42560 1 0 $X=19730 $Y=37440
X9923 3 1 DECAP7JI3V $T=20160 51520 0 0 $X=19730 $Y=50880
X9924 3 1 DECAP7JI3V $T=20160 78400 1 0 $X=19730 $Y=73280
X9925 3 1 DECAP7JI3V $T=20160 78400 0 0 $X=19730 $Y=77760
X9926 3 1 DECAP7JI3V $T=20160 105280 1 0 $X=19730 $Y=100160
X9927 3 1 DECAP7JI3V $T=20160 105280 0 0 $X=19730 $Y=104640
X9928 3 1 DECAP7JI3V $T=20160 114240 1 0 $X=19730 $Y=109120
X9929 3 1 DECAP7JI3V $T=20160 114240 0 0 $X=19730 $Y=113600
X9930 3 1 DECAP7JI3V $T=20160 123200 0 0 $X=19730 $Y=122560
X9931 3 1 DECAP7JI3V $T=20160 141120 1 0 $X=19730 $Y=136000
X9932 3 1 DECAP7JI3V $T=20160 141120 0 0 $X=19730 $Y=140480
X9933 3 1 DECAP7JI3V $T=20160 159040 0 0 $X=19730 $Y=158400
X9934 3 1 DECAP7JI3V $T=20160 185920 1 0 $X=19730 $Y=180800
X9935 3 1 DECAP7JI3V $T=20160 185920 0 0 $X=19730 $Y=185280
X9936 3 1 DECAP7JI3V $T=20160 194880 0 0 $X=19730 $Y=194240
X9937 3 1 DECAP7JI3V $T=20160 203840 1 0 $X=19730 $Y=198720
X9938 3 1 DECAP7JI3V $T=24080 78400 0 0 $X=23650 $Y=77760
X9939 3 1 DECAP7JI3V $T=24080 159040 0 0 $X=23650 $Y=158400
X9940 3 1 DECAP7JI3V $T=24080 203840 1 0 $X=23650 $Y=198720
X9941 3 1 DECAP7JI3V $T=28000 203840 1 0 $X=27570 $Y=198720
X9942 3 1 DECAP7JI3V $T=31920 203840 1 0 $X=31490 $Y=198720
X9943 3 1 DECAP7JI3V $T=34160 24640 0 0 $X=33730 $Y=24000
X9944 3 1 DECAP7JI3V $T=34160 168000 1 0 $X=33730 $Y=162880
X9945 3 1 DECAP7JI3V $T=34720 114240 0 0 $X=34290 $Y=113600
X9946 3 1 DECAP7JI3V $T=34720 123200 1 0 $X=34290 $Y=118080
X9947 3 1 DECAP7JI3V $T=38080 24640 0 0 $X=37650 $Y=24000
X9948 3 1 DECAP7JI3V $T=38080 168000 1 0 $X=37650 $Y=162880
X9949 3 1 DECAP7JI3V $T=38640 123200 1 0 $X=38210 $Y=118080
X9950 3 1 DECAP7JI3V $T=42000 24640 0 0 $X=41570 $Y=24000
X9951 3 1 DECAP7JI3V $T=42000 168000 1 0 $X=41570 $Y=162880
X9952 3 1 DECAP7JI3V $T=43120 42560 0 0 $X=42690 $Y=41920
X9953 3 1 DECAP7JI3V $T=43120 78400 0 0 $X=42690 $Y=77760
X9954 3 1 DECAP7JI3V $T=43680 123200 1 0 $X=43250 $Y=118080
X9955 3 1 DECAP7JI3V $T=45920 24640 0 0 $X=45490 $Y=24000
X9956 3 1 DECAP7JI3V $T=49280 159040 0 0 $X=48850 $Y=158400
X9957 3 1 DECAP7JI3V $T=53760 24640 1 0 $X=53330 $Y=19520
X9958 3 1 DECAP7JI3V $T=53760 221760 1 0 $X=53330 $Y=216640
X9959 3 1 DECAP7JI3V $T=57680 24640 1 0 $X=57250 $Y=19520
X9960 3 1 DECAP7JI3V $T=57680 221760 1 0 $X=57250 $Y=216640
X9961 3 1 DECAP7JI3V $T=62720 150080 0 0 $X=62290 $Y=149440
X9962 3 1 DECAP7JI3V $T=64400 176960 1 0 $X=63970 $Y=171840
X9963 3 1 DECAP7JI3V $T=69440 78400 1 0 $X=69010 $Y=73280
X9964 3 1 DECAP7JI3V $T=77280 60480 0 0 $X=76850 $Y=59840
X9965 3 1 DECAP7JI3V $T=92960 33600 0 180 $X=88610 $Y=28480
X9966 3 1 DECAP7JI3V $T=94640 87360 1 0 $X=94210 $Y=82240
X9967 3 1 DECAP7JI3V $T=101360 60480 1 0 $X=100930 $Y=55360
X9968 3 1 DECAP7JI3V $T=101360 60480 0 0 $X=100930 $Y=59840
X9969 3 1 DECAP7JI3V $T=101360 69440 1 0 $X=100930 $Y=64320
X9970 3 1 DECAP7JI3V $T=101360 69440 0 0 $X=100930 $Y=68800
X9971 3 1 DECAP7JI3V $T=101360 78400 1 0 $X=100930 $Y=73280
X9972 3 1 DECAP7JI3V $T=101360 168000 0 0 $X=100930 $Y=167360
X9973 3 1 DECAP7JI3V $T=103040 105280 0 0 $X=102610 $Y=104640
X9974 3 1 DECAP7JI3V $T=105280 24640 1 0 $X=104850 $Y=19520
X9975 3 1 DECAP7JI3V $T=105280 42560 0 0 $X=104850 $Y=41920
X9976 3 1 DECAP7JI3V $T=105280 51520 0 0 $X=104850 $Y=50880
X9977 3 1 DECAP7JI3V $T=105280 60480 1 0 $X=104850 $Y=55360
X9978 3 1 DECAP7JI3V $T=105280 60480 0 0 $X=104850 $Y=59840
X9979 3 1 DECAP7JI3V $T=105280 69440 1 0 $X=104850 $Y=64320
X9980 3 1 DECAP7JI3V $T=105280 69440 0 0 $X=104850 $Y=68800
X9981 3 1 DECAP7JI3V $T=105280 78400 1 0 $X=104850 $Y=73280
X9982 3 1 DECAP7JI3V $T=105280 87360 1 0 $X=104850 $Y=82240
X9983 3 1 DECAP7JI3V $T=105280 132160 1 0 $X=104850 $Y=127040
X9984 3 1 DECAP7JI3V $T=105280 132160 0 0 $X=104850 $Y=131520
X9985 3 1 DECAP7JI3V $T=105280 141120 1 0 $X=104850 $Y=136000
X9986 3 1 DECAP7JI3V $T=105280 141120 0 0 $X=104850 $Y=140480
X9987 3 1 DECAP7JI3V $T=105280 150080 1 0 $X=104850 $Y=144960
X9988 3 1 DECAP7JI3V $T=105280 194880 0 0 $X=104850 $Y=194240
X9989 3 1 DECAP7JI3V $T=106400 176960 1 0 $X=105970 $Y=171840
X9990 3 1 DECAP7JI3V $T=106960 105280 0 0 $X=106530 $Y=104640
X9991 3 1 DECAP7JI3V $T=109200 24640 1 0 $X=108770 $Y=19520
X9992 3 1 DECAP7JI3V $T=109200 60480 1 0 $X=108770 $Y=55360
X9993 3 1 DECAP7JI3V $T=109200 60480 0 0 $X=108770 $Y=59840
X9994 3 1 DECAP7JI3V $T=109200 69440 1 0 $X=108770 $Y=64320
X9995 3 1 DECAP7JI3V $T=109200 69440 0 0 $X=108770 $Y=68800
X9996 3 1 DECAP7JI3V $T=109200 78400 1 0 $X=108770 $Y=73280
X9997 3 1 DECAP7JI3V $T=109200 87360 1 0 $X=108770 $Y=82240
X9998 3 1 DECAP7JI3V $T=109200 132160 1 0 $X=108770 $Y=127040
X9999 3 1 DECAP7JI3V $T=109200 132160 0 0 $X=108770 $Y=131520
X10000 3 1 DECAP7JI3V $T=109200 141120 1 0 $X=108770 $Y=136000
X10001 3 1 DECAP7JI3V $T=109200 141120 0 0 $X=108770 $Y=140480
X10002 3 1 DECAP7JI3V $T=109200 150080 1 0 $X=108770 $Y=144960
X10003 3 1 DECAP7JI3V $T=109200 159040 0 0 $X=108770 $Y=158400
X10004 3 1 DECAP7JI3V $T=109200 194880 0 0 $X=108770 $Y=194240
X10005 3 1 DECAP7JI3V $T=110320 176960 1 0 $X=109890 $Y=171840
X10006 3 1 DECAP7JI3V $T=114240 176960 1 0 $X=113810 $Y=171840
X10007 3 1 DECAP7JI3V $T=118720 78400 1 0 $X=118290 $Y=73280
X10008 3 1 DECAP7JI3V $T=118720 150080 0 0 $X=118290 $Y=149440
X10009 3 1 DECAP7JI3V $T=118720 212800 1 0 $X=118290 $Y=207680
X10010 3 1 DECAP7JI3V $T=118720 221760 1 0 $X=118290 $Y=216640
X10011 3 1 DECAP7JI3V $T=123200 168000 1 0 $X=122770 $Y=162880
X10012 3 1 DECAP7JI3V $T=123200 168000 0 0 $X=122770 $Y=167360
X10013 3 1 DECAP7JI3V $T=127120 212800 1 180 $X=122770 $Y=212160
X10014 3 1 DECAP7JI3V $T=127120 212800 0 0 $X=126690 $Y=212160
X10015 3 1 DECAP7JI3V $T=132720 33600 1 180 $X=128370 $Y=32960
X10016 3 1 DECAP7JI3V $T=131040 212800 0 0 $X=130610 $Y=212160
X10017 3 1 DECAP7JI3V $T=132720 185920 1 0 $X=132290 $Y=180800
X10018 3 1 DECAP7JI3V $T=133280 132160 0 0 $X=132850 $Y=131520
X10019 3 1 DECAP7JI3V $T=134960 212800 0 0 $X=134530 $Y=212160
X10020 3 1 DECAP7JI3V $T=149520 78400 0 0 $X=149090 $Y=77760
X10021 3 1 DECAP7JI3V $T=153440 78400 0 0 $X=153010 $Y=77760
X10022 3 1 DECAP7JI3V $T=154000 96320 1 0 $X=153570 $Y=91200
X10023 3 1 DECAP7JI3V $T=157360 78400 0 0 $X=156930 $Y=77760
X10024 3 1 DECAP7JI3V $T=157920 96320 1 0 $X=157490 $Y=91200
X10025 3 1 DECAP7JI3V $T=159040 123200 1 0 $X=158610 $Y=118080
X10026 3 1 DECAP7JI3V $T=161280 78400 0 0 $X=160850 $Y=77760
X10027 3 1 DECAP7JI3V $T=161840 96320 1 0 $X=161410 $Y=91200
X10028 3 1 DECAP7JI3V $T=162960 123200 1 0 $X=162530 $Y=118080
X10029 3 1 DECAP7JI3V $T=167440 105280 1 0 $X=167010 $Y=100160
X10030 3 1 DECAP7JI3V $T=174160 33600 0 0 $X=173730 $Y=32960
X10031 3 1 DECAP7JI3V $T=175840 141120 0 0 $X=175410 $Y=140480
X10032 3 1 DECAP7JI3V $T=179200 132160 1 0 $X=178770 $Y=127040
X10033 3 1 DECAP7JI3V $T=180320 105280 0 0 $X=179890 $Y=104640
X10034 3 1 DECAP7JI3V $T=182560 78400 1 0 $X=182130 $Y=73280
X10035 3 1 DECAP7JI3V $T=184240 33600 1 0 $X=183810 $Y=28480
X10036 3 1 DECAP7JI3V $T=184240 60480 1 0 $X=183810 $Y=55360
X10037 3 1 DECAP7JI3V $T=184240 105280 0 0 $X=183810 $Y=104640
X10038 3 1 DECAP7JI3V $T=185920 87360 1 0 $X=185490 $Y=82240
X10039 3 1 DECAP7JI3V $T=185920 132160 1 0 $X=185490 $Y=127040
X10040 3 1 DECAP7JI3V $T=190400 78400 0 180 $X=186050 $Y=73280
X10041 3 1 DECAP7JI3V $T=189840 87360 1 0 $X=189410 $Y=82240
X10042 3 1 DECAP7JI3V $T=194880 60480 0 0 $X=194450 $Y=59840
X10043 3 1 DECAP7JI3V $T=203280 123200 0 0 $X=202850 $Y=122560
X10044 3 1 DECAP7JI3V $T=203280 132160 0 0 $X=202850 $Y=131520
X10045 3 1 DECAP7JI3V $T=206080 168000 1 0 $X=205650 $Y=162880
X10046 3 1 DECAP7JI3V $T=206080 168000 0 0 $X=205650 $Y=167360
X10047 3 1 DECAP7JI3V $T=206080 176960 1 0 $X=205650 $Y=171840
X10048 3 1 DECAP7JI3V $T=207200 123200 0 0 $X=206770 $Y=122560
X10049 3 1 DECAP7JI3V $T=207200 132160 0 0 $X=206770 $Y=131520
X10050 3 1 DECAP7JI3V $T=207200 150080 0 0 $X=206770 $Y=149440
X10051 3 1 DECAP7JI3V $T=208320 105280 0 0 $X=207890 $Y=104640
X10052 3 1 DECAP7JI3V $T=210000 168000 1 0 $X=209570 $Y=162880
X10053 3 1 DECAP7JI3V $T=210000 168000 0 0 $X=209570 $Y=167360
X10054 3 1 DECAP7JI3V $T=210000 176960 1 0 $X=209570 $Y=171840
X10055 3 1 DECAP7JI3V $T=211120 96320 0 0 $X=210690 $Y=95680
X10056 3 1 DECAP7JI3V $T=211120 123200 0 0 $X=210690 $Y=122560
X10057 3 1 DECAP7JI3V $T=211120 132160 1 0 $X=210690 $Y=127040
X10058 3 1 DECAP7JI3V $T=211120 132160 0 0 $X=210690 $Y=131520
X10059 3 1 DECAP7JI3V $T=211120 150080 0 0 $X=210690 $Y=149440
X10060 3 1 DECAP7JI3V $T=212240 105280 0 0 $X=211810 $Y=104640
X10061 3 1 DECAP7JI3V $T=213920 114240 0 0 $X=213490 $Y=113600
X10062 3 1 DECAP7JI3V $T=215040 96320 0 0 $X=214610 $Y=95680
X10063 3 1 DECAP7JI3V $T=215040 123200 0 0 $X=214610 $Y=122560
X10064 3 1 DECAP7JI3V $T=215040 132160 1 0 $X=214610 $Y=127040
X10065 3 1 DECAP7JI3V $T=215040 132160 0 0 $X=214610 $Y=131520
X10066 3 1 DECAP7JI3V $T=215040 141120 1 0 $X=214610 $Y=136000
X10067 3 1 DECAP7JI3V $T=215040 150080 0 0 $X=214610 $Y=149440
X10068 3 1 DECAP7JI3V $T=215040 159040 0 0 $X=214610 $Y=158400
X10069 3 1 DECAP7JI3V $T=215040 176960 0 0 $X=214610 $Y=176320
X10070 3 1 DECAP7JI3V $T=218960 141120 1 0 $X=218530 $Y=136000
X10071 3 1 DECAP7JI3V $T=236320 42560 1 0 $X=235890 $Y=37440
X10072 3 1 DECAP7JI3V $T=243600 87360 1 0 $X=243170 $Y=82240
X10073 3 1 DECAP7JI3V $T=254800 168000 1 180 $X=250450 $Y=167360
X10074 3 1 DECAP7JI3V $T=253680 141120 1 0 $X=253250 $Y=136000
X10075 3 1 DECAP7JI3V $T=261520 141120 0 180 $X=257170 $Y=136000
X10076 3 1 DECAP7JI3V $T=260400 87360 0 0 $X=259970 $Y=86720
X10077 3 1 DECAP7JI3V $T=260400 123200 1 0 $X=259970 $Y=118080
X10078 3 1 DECAP7JI3V $T=260400 123200 0 0 $X=259970 $Y=122560
X10079 3 1 DECAP7JI3V $T=260960 132160 1 0 $X=260530 $Y=127040
X10080 3 1 DECAP7JI3V $T=264320 87360 0 0 $X=263890 $Y=86720
X10081 3 1 DECAP7JI3V $T=268240 87360 0 0 $X=267810 $Y=86720
X10082 3 1 DECAP7JI3V $T=277200 176960 0 0 $X=276770 $Y=176320
X10083 3 1 DECAP7JI3V $T=278880 78400 0 0 $X=278450 $Y=77760
X10084 3 1 DECAP7JI3V $T=282240 105280 1 0 $X=281810 $Y=100160
X10085 3 1 DECAP7JI3V $T=282240 114240 1 0 $X=281810 $Y=109120
X10086 3 1 DECAP7JI3V $T=282800 78400 0 0 $X=282370 $Y=77760
X10087 3 1 DECAP7JI3V $T=284480 123200 0 0 $X=284050 $Y=122560
X10088 3 1 DECAP7JI3V $T=285040 132160 0 0 $X=284610 $Y=131520
X10089 3 1 DECAP7JI3V $T=286160 105280 1 0 $X=285730 $Y=100160
X10090 3 1 DECAP7JI3V $T=290080 105280 1 0 $X=289650 $Y=100160
X10091 3 1 DECAP7JI3V $T=290640 96320 1 0 $X=290210 $Y=91200
X10092 3 1 DECAP7JI3V $T=293440 87360 0 0 $X=293010 $Y=86720
X10093 3 1 DECAP7JI3V $T=297360 87360 0 0 $X=296930 $Y=86720
X10094 3 1 DECAP7JI3V $T=305760 42560 0 0 $X=305330 $Y=41920
X10095 3 1 DECAP7JI3V $T=306880 42560 1 0 $X=306450 $Y=37440
X10096 3 1 DECAP7JI3V $T=307440 150080 1 0 $X=307010 $Y=144960
X10097 3 1 DECAP7JI3V $T=309120 78400 1 0 $X=308690 $Y=73280
X10098 3 1 DECAP7JI3V $T=309120 96320 0 0 $X=308690 $Y=95680
X10099 3 1 DECAP7JI3V $T=309120 105280 1 0 $X=308690 $Y=100160
X10100 3 1 DECAP7JI3V $T=309120 114240 1 0 $X=308690 $Y=109120
X10101 3 1 DECAP7JI3V $T=309120 141120 0 0 $X=308690 $Y=140480
X10102 3 1 DECAP7JI3V $T=313040 78400 1 0 $X=312610 $Y=73280
X10103 3 1 DECAP7JI3V $T=313040 96320 0 0 $X=312610 $Y=95680
X10104 3 1 DECAP7JI3V $T=313040 105280 1 0 $X=312610 $Y=100160
X10105 3 1 DECAP7JI3V $T=313040 114240 1 0 $X=312610 $Y=109120
X10106 3 1 DECAP7JI3V $T=313040 141120 0 0 $X=312610 $Y=140480
X10107 3 1 DECAP7JI3V $T=315840 141120 1 0 $X=315410 $Y=136000
X10108 3 1 DECAP7JI3V $T=315840 159040 0 0 $X=315410 $Y=158400
X10109 3 1 DECAP7JI3V $T=315840 168000 1 0 $X=315410 $Y=162880
X10110 3 1 DECAP7JI3V $T=316960 78400 1 0 $X=316530 $Y=73280
X10111 3 1 DECAP7JI3V $T=316960 123200 1 0 $X=316530 $Y=118080
X10112 3 1 DECAP7JI3V $T=316960 132160 1 0 $X=316530 $Y=127040
X10113 3 1 DECAP7JI3V $T=316960 150080 1 0 $X=316530 $Y=144960
X10114 3 1 DECAP7JI3V $T=318080 87360 0 0 $X=317650 $Y=86720
X10115 3 1 DECAP7JI3V $T=318080 123200 0 0 $X=317650 $Y=122560
X10116 3 1 DECAP7JI3V $T=319200 42560 0 0 $X=318770 $Y=41920
X10117 3 1 DECAP7JI3V $T=320880 69440 0 0 $X=320450 $Y=68800
X10118 3 1 DECAP7JI3V $T=320880 78400 1 0 $X=320450 $Y=73280
X10119 3 1 DECAP7JI3V $T=320880 87360 1 0 $X=320450 $Y=82240
X10120 3 1 DECAP7JI3V $T=320880 123200 1 0 $X=320450 $Y=118080
X10121 3 1 DECAP7JI3V $T=320880 132160 1 0 $X=320450 $Y=127040
X10122 3 1 DECAP7JI3V $T=320880 150080 1 0 $X=320450 $Y=144960
X10123 3 1 DECAP7JI3V $T=322000 212800 1 0 $X=321570 $Y=207680
X10124 3 1 DECAP7JI3V $T=329840 132160 0 0 $X=329410 $Y=131520
X10125 3 1 DECAP7JI3V $T=330400 78400 0 0 $X=329970 $Y=77760
X10126 3 1 DECAP7JI3V $T=330400 105280 0 0 $X=329970 $Y=104640
X10127 3 1 DECAP7JI3V $T=334320 78400 0 0 $X=333890 $Y=77760
X10128 3 1 DECAP7JI3V $T=344960 114240 0 0 $X=344530 $Y=113600
X10129 3 1 DECAP7JI3V $T=348880 114240 0 0 $X=348450 $Y=113600
X10130 3 1 DECAP7JI3V $T=352800 114240 0 0 $X=352370 $Y=113600
X10131 3 1 DECAP7JI3V $T=352800 141120 0 0 $X=352370 $Y=140480
X10132 3 1 DECAP7JI3V $T=356720 114240 1 0 $X=356290 $Y=109120
X10133 3 1 DECAP7JI3V $T=356720 114240 0 0 $X=356290 $Y=113600
X10134 3 1 DECAP7JI3V $T=356720 141120 0 0 $X=356290 $Y=140480
X10135 3 1 DECAP7JI3V $T=357280 42560 0 0 $X=356850 $Y=41920
X10136 3 1 DECAP7JI3V $T=357280 51520 1 0 $X=356850 $Y=46400
X10137 3 1 DECAP7JI3V $T=358400 96320 1 0 $X=357970 $Y=91200
X10138 3 1 DECAP7JI3V $T=358960 60480 1 0 $X=358530 $Y=55360
X10139 3 1 DECAP7JI3V $T=359520 78400 0 0 $X=359090 $Y=77760
X10140 3 1 DECAP7JI3V $T=360080 69440 0 0 $X=359650 $Y=68800
X10141 3 1 DECAP7JI3V $T=406560 78400 0 0 $X=406130 $Y=77760
X10142 3 1 DECAP7JI3V $T=406560 87360 0 0 $X=406130 $Y=86720
X10143 3 1 DECAP7JI3V $T=406560 96320 1 0 $X=406130 $Y=91200
X10144 3 1 DECAP7JI3V $T=406560 150080 0 0 $X=406130 $Y=149440
X10145 3 1 DECAP7JI3V $T=409360 78400 1 0 $X=408930 $Y=73280
X10146 3 1 DECAP7JI3V $T=409360 87360 1 0 $X=408930 $Y=82240
X10147 3 1 DECAP7JI3V $T=409360 150080 1 0 $X=408930 $Y=144960
X10148 3 1 DECAP7JI3V $T=409360 203840 1 0 $X=408930 $Y=198720
X10149 3 1 DECAP7JI3V $T=409360 212800 1 0 $X=408930 $Y=207680
X10150 3 1 DECAP7JI3V $T=410480 69440 1 0 $X=410050 $Y=64320
X10151 3 1 DECAP7JI3V $T=410480 78400 0 0 $X=410050 $Y=77760
X10152 3 1 DECAP7JI3V $T=410480 87360 0 0 $X=410050 $Y=86720
X10153 3 1 DECAP7JI3V $T=410480 96320 1 0 $X=410050 $Y=91200
X10154 3 1 DECAP7JI3V $T=410480 150080 0 0 $X=410050 $Y=149440
X10155 3 1 DECAP7JI3V $T=410480 185920 1 0 $X=410050 $Y=180800
X10156 3 1 DECAP7JI3V $T=413280 33600 0 0 $X=412850 $Y=32960
X10157 3 1 DECAP7JI3V $T=413280 78400 1 0 $X=412850 $Y=73280
X10158 3 1 DECAP7JI3V $T=413280 87360 1 0 $X=412850 $Y=82240
X10159 3 1 DECAP7JI3V $T=413280 150080 1 0 $X=412850 $Y=144960
X10160 3 1 DECAP7JI3V $T=413280 194880 0 0 $X=412850 $Y=194240
X10161 3 1 DECAP7JI3V $T=413280 203840 1 0 $X=412850 $Y=198720
X10162 3 1 DECAP7JI3V $T=413280 203840 0 0 $X=412850 $Y=203200
X10163 3 1 DECAP7JI3V $T=413280 212800 1 0 $X=412850 $Y=207680
X10164 3 1 DECAP7JI3V $T=414400 69440 1 0 $X=413970 $Y=64320
X10165 3 1 DECAP7JI3V $T=414400 78400 0 0 $X=413970 $Y=77760
X10166 3 1 DECAP7JI3V $T=414400 87360 0 0 $X=413970 $Y=86720
X10167 3 1 DECAP7JI3V $T=414400 96320 1 0 $X=413970 $Y=91200
X10168 3 1 DECAP7JI3V $T=414400 105280 0 0 $X=413970 $Y=104640
X10169 3 1 DECAP7JI3V $T=414400 123200 1 0 $X=413970 $Y=118080
X10170 3 1 DECAP7JI3V $T=414400 150080 0 0 $X=413970 $Y=149440
X10171 3 1 DECAP7JI3V $T=414400 176960 0 0 $X=413970 $Y=176320
X10172 3 1 DECAP7JI3V $T=414400 185920 1 0 $X=413970 $Y=180800
X10173 3 1 DECAP7JI3V $T=414400 194880 1 0 $X=413970 $Y=189760
X10174 3 1 DECAP7JI3V $T=414400 212800 0 0 $X=413970 $Y=212160
X10175 3 1 DECAP7JI3V $T=417200 33600 1 0 $X=416770 $Y=28480
X10176 3 1 DECAP7JI3V $T=417200 33600 0 0 $X=416770 $Y=32960
X10177 3 1 DECAP7JI3V $T=417200 78400 1 0 $X=416770 $Y=73280
X10178 3 1 DECAP7JI3V $T=417200 87360 1 0 $X=416770 $Y=82240
X10179 3 1 DECAP7JI3V $T=417200 114240 1 0 $X=416770 $Y=109120
X10180 3 1 DECAP7JI3V $T=417200 123200 0 0 $X=416770 $Y=122560
X10181 3 1 DECAP7JI3V $T=417200 141120 0 0 $X=416770 $Y=140480
X10182 3 1 DECAP7JI3V $T=417200 150080 1 0 $X=416770 $Y=144960
X10183 3 1 DECAP7JI3V $T=417200 194880 0 0 $X=416770 $Y=194240
X10184 3 1 DECAP7JI3V $T=417200 203840 1 0 $X=416770 $Y=198720
X10185 3 1 DECAP7JI3V $T=417200 203840 0 0 $X=416770 $Y=203200
X10186 3 1 DECAP7JI3V $T=417200 212800 1 0 $X=416770 $Y=207680
X10187 3 1 DECAP7JI3V $T=418320 69440 1 0 $X=417890 $Y=64320
X10188 3 1 DECAP7JI3V $T=418320 78400 0 0 $X=417890 $Y=77760
X10189 3 1 DECAP7JI3V $T=418320 87360 0 0 $X=417890 $Y=86720
X10190 3 1 DECAP7JI3V $T=418320 96320 1 0 $X=417890 $Y=91200
X10191 3 1 DECAP7JI3V $T=418320 96320 0 0 $X=417890 $Y=95680
X10192 3 1 DECAP7JI3V $T=418320 105280 1 0 $X=417890 $Y=100160
X10193 3 1 DECAP7JI3V $T=418320 105280 0 0 $X=417890 $Y=104640
X10194 3 1 DECAP7JI3V $T=418320 114240 0 0 $X=417890 $Y=113600
X10195 3 1 DECAP7JI3V $T=418320 123200 1 0 $X=417890 $Y=118080
X10196 3 1 DECAP7JI3V $T=418320 132160 0 0 $X=417890 $Y=131520
X10197 3 1 DECAP7JI3V $T=418320 141120 1 0 $X=417890 $Y=136000
X10198 3 1 DECAP7JI3V $T=418320 150080 0 0 $X=417890 $Y=149440
X10199 3 1 DECAP7JI3V $T=418320 176960 0 0 $X=417890 $Y=176320
X10200 3 1 DECAP7JI3V $T=418320 185920 1 0 $X=417890 $Y=180800
X10201 3 1 DECAP7JI3V $T=418320 194880 1 0 $X=417890 $Y=189760
X10202 3 1 DECAP7JI3V $T=418320 212800 0 0 $X=417890 $Y=212160
X10203 3 1 DECAP7JI3V $T=421120 33600 1 0 $X=420690 $Y=28480
X10204 3 1 DECAP7JI3V $T=421120 33600 0 0 $X=420690 $Y=32960
X10205 3 1 DECAP7JI3V $T=421120 42560 1 0 $X=420690 $Y=37440
X10206 3 1 DECAP7JI3V $T=421120 42560 0 0 $X=420690 $Y=41920
X10207 3 1 DECAP7JI3V $T=421120 51520 1 0 $X=420690 $Y=46400
X10208 3 1 DECAP7JI3V $T=421120 51520 0 0 $X=420690 $Y=50880
X10209 3 1 DECAP7JI3V $T=421120 60480 1 0 $X=420690 $Y=55360
X10210 3 1 DECAP7JI3V $T=421120 60480 0 0 $X=420690 $Y=59840
X10211 3 1 DECAP7JI3V $T=421120 69440 0 0 $X=420690 $Y=68800
X10212 3 1 DECAP7JI3V $T=421120 78400 1 0 $X=420690 $Y=73280
X10213 3 1 DECAP7JI3V $T=421120 87360 1 0 $X=420690 $Y=82240
X10214 3 1 DECAP7JI3V $T=421120 114240 1 0 $X=420690 $Y=109120
X10215 3 1 DECAP7JI3V $T=421120 123200 0 0 $X=420690 $Y=122560
X10216 3 1 DECAP7JI3V $T=421120 132160 1 0 $X=420690 $Y=127040
X10217 3 1 DECAP7JI3V $T=421120 141120 0 0 $X=420690 $Y=140480
X10218 3 1 DECAP7JI3V $T=421120 150080 1 0 $X=420690 $Y=144960
X10219 3 1 DECAP7JI3V $T=421120 159040 0 0 $X=420690 $Y=158400
X10220 3 1 DECAP7JI3V $T=421120 168000 1 0 $X=420690 $Y=162880
X10221 3 1 DECAP7JI3V $T=421120 168000 0 0 $X=420690 $Y=167360
X10222 3 1 DECAP7JI3V $T=421120 176960 1 0 $X=420690 $Y=171840
X10223 3 1 DECAP7JI3V $T=421120 194880 0 0 $X=420690 $Y=194240
X10224 3 1 DECAP7JI3V $T=421120 203840 1 0 $X=420690 $Y=198720
X10225 3 1 DECAP7JI3V $T=421120 203840 0 0 $X=420690 $Y=203200
X10226 3 1 DECAP7JI3V $T=421120 212800 1 0 $X=420690 $Y=207680
X10227 3 1 DECAP5JI3V $T=20160 42560 0 0 $X=19730 $Y=41920
X10228 3 1 DECAP5JI3V $T=20160 51520 1 0 $X=19730 $Y=46400
X10229 3 1 DECAP5JI3V $T=20160 96320 0 0 $X=19730 $Y=95680
X10230 3 1 DECAP5JI3V $T=20160 132160 1 0 $X=19730 $Y=127040
X10231 3 1 DECAP5JI3V $T=20160 159040 1 0 $X=19730 $Y=153920
X10232 3 1 DECAP5JI3V $T=20160 176960 1 0 $X=19730 $Y=171840
X10233 3 1 DECAP5JI3V $T=30800 78400 1 180 $X=27570 $Y=77760
X10234 3 1 DECAP5JI3V $T=28560 203840 0 0 $X=28130 $Y=203200
X10235 3 1 DECAP5JI3V $T=34720 132160 1 0 $X=34290 $Y=127040
X10236 3 1 DECAP5JI3V $T=38640 203840 0 180 $X=35410 $Y=198720
X10237 3 1 DECAP5JI3V $T=39200 123200 0 0 $X=38770 $Y=122560
X10238 3 1 DECAP5JI3V $T=40880 96320 1 0 $X=40450 $Y=91200
X10239 3 1 DECAP5JI3V $T=42560 212800 0 0 $X=42130 $Y=212160
X10240 3 1 DECAP5JI3V $T=49840 24640 0 0 $X=49410 $Y=24000
X10241 3 1 DECAP5JI3V $T=57120 51520 0 0 $X=56690 $Y=50880
X10242 3 1 DECAP5JI3V $T=59360 60480 0 0 $X=58930 $Y=59840
X10243 3 1 DECAP5JI3V $T=59360 87360 1 0 $X=58930 $Y=82240
X10244 3 1 DECAP5JI3V $T=61040 33600 1 0 $X=60610 $Y=28480
X10245 3 1 DECAP5JI3V $T=66640 150080 0 0 $X=66210 $Y=149440
X10246 3 1 DECAP5JI3V $T=76720 60480 1 0 $X=76290 $Y=55360
X10247 3 1 DECAP5JI3V $T=78400 33600 0 0 $X=77970 $Y=32960
X10248 3 1 DECAP5JI3V $T=84000 105280 0 0 $X=83570 $Y=104640
X10249 3 1 DECAP5JI3V $T=105280 105280 1 0 $X=104850 $Y=100160
X10250 3 1 DECAP5JI3V $T=105280 168000 0 0 $X=104850 $Y=167360
X10251 3 1 DECAP5JI3V $T=105280 176960 0 0 $X=104850 $Y=176320
X10252 3 1 DECAP5JI3V $T=105280 212800 0 0 $X=104850 $Y=212160
X10253 3 1 DECAP5JI3V $T=108640 150080 0 0 $X=108210 $Y=149440
X10254 3 1 DECAP5JI3V $T=108640 159040 1 0 $X=108210 $Y=153920
X10255 3 1 DECAP5JI3V $T=110320 96320 0 0 $X=109890 $Y=95680
X10256 3 1 DECAP5JI3V $T=110320 203840 1 0 $X=109890 $Y=198720
X10257 3 1 DECAP5JI3V $T=113120 123200 1 0 $X=112690 $Y=118080
X10258 3 1 DECAP5JI3V $T=113120 159040 0 0 $X=112690 $Y=158400
X10259 3 1 DECAP5JI3V $T=122640 78400 1 0 $X=122210 $Y=73280
X10260 3 1 DECAP5JI3V $T=122640 150080 0 0 $X=122210 $Y=149440
X10261 3 1 DECAP5JI3V $T=133280 114240 0 0 $X=132850 $Y=113600
X10262 3 1 DECAP5JI3V $T=143360 212800 1 0 $X=142930 $Y=207680
X10263 3 1 DECAP5JI3V $T=156240 132160 1 0 $X=155810 $Y=127040
X10264 3 1 DECAP5JI3V $T=164080 87360 1 0 $X=163650 $Y=82240
X10265 3 1 DECAP5JI3V $T=166880 123200 1 0 $X=166450 $Y=118080
X10266 3 1 DECAP5JI3V $T=168560 96320 0 0 $X=168130 $Y=95680
X10267 3 1 DECAP5JI3V $T=179760 141120 0 0 $X=179330 $Y=140480
X10268 3 1 DECAP5JI3V $T=188160 150080 1 0 $X=187730 $Y=144960
X10269 3 1 DECAP5JI3V $T=190960 168000 1 180 $X=187730 $Y=167360
X10270 3 1 DECAP5JI3V $T=188160 176960 1 0 $X=187730 $Y=171840
X10271 3 1 DECAP5JI3V $T=211120 185920 1 0 $X=210690 $Y=180800
X10272 3 1 DECAP5JI3V $T=211120 212800 1 0 $X=210690 $Y=207680
X10273 3 1 DECAP5JI3V $T=211680 42560 0 0 $X=211250 $Y=41920
X10274 3 1 DECAP5JI3V $T=211680 51520 1 0 $X=211250 $Y=46400
X10275 3 1 DECAP5JI3V $T=211680 60480 1 0 $X=211250 $Y=55360
X10276 3 1 DECAP5JI3V $T=211680 69440 0 0 $X=211250 $Y=68800
X10277 3 1 DECAP5JI3V $T=211680 78400 0 0 $X=211250 $Y=77760
X10278 3 1 DECAP5JI3V $T=214480 87360 0 0 $X=214050 $Y=86720
X10279 3 1 DECAP5JI3V $T=214480 150080 1 0 $X=214050 $Y=144960
X10280 3 1 DECAP5JI3V $T=215040 212800 0 0 $X=214610 $Y=212160
X10281 3 1 DECAP5JI3V $T=216160 96320 1 0 $X=215730 $Y=91200
X10282 3 1 DECAP5JI3V $T=216160 105280 0 0 $X=215730 $Y=104640
X10283 3 1 DECAP5JI3V $T=229600 42560 0 0 $X=229170 $Y=41920
X10284 3 1 DECAP5JI3V $T=232400 51520 0 180 $X=229170 $Y=46400
X10285 3 1 DECAP5JI3V $T=229600 60480 1 0 $X=229170 $Y=55360
X10286 3 1 DECAP5JI3V $T=230720 168000 1 0 $X=230290 $Y=162880
X10287 3 1 DECAP5JI3V $T=239120 141120 0 0 $X=238690 $Y=140480
X10288 3 1 DECAP5JI3V $T=247520 51520 0 0 $X=247090 $Y=50880
X10289 3 1 DECAP5JI3V $T=250320 60480 0 180 $X=247090 $Y=55360
X10290 3 1 DECAP5JI3V $T=261520 141120 1 0 $X=261090 $Y=136000
X10291 3 1 DECAP5JI3V $T=267680 96320 1 0 $X=267250 $Y=91200
X10292 3 1 DECAP5JI3V $T=269360 78400 1 0 $X=268930 $Y=73280
X10293 3 1 DECAP5JI3V $T=274400 114240 0 0 $X=273970 $Y=113600
X10294 3 1 DECAP5JI3V $T=284480 105280 0 0 $X=284050 $Y=104640
X10295 3 1 DECAP5JI3V $T=285600 123200 1 0 $X=285170 $Y=118080
X10296 3 1 DECAP5JI3V $T=286160 114240 1 0 $X=285730 $Y=109120
X10297 3 1 DECAP5JI3V $T=286160 141120 1 0 $X=285730 $Y=136000
X10298 3 1 DECAP5JI3V $T=289520 78400 1 180 $X=286290 $Y=77760
X10299 3 1 DECAP5JI3V $T=291200 96320 0 0 $X=290770 $Y=95680
X10300 3 1 DECAP5JI3V $T=301280 87360 0 0 $X=300850 $Y=86720
X10301 3 1 DECAP5JI3V $T=309120 194880 1 0 $X=308690 $Y=189760
X10302 3 1 DECAP5JI3V $T=316960 51520 0 0 $X=316530 $Y=50880
X10303 3 1 DECAP5JI3V $T=316960 60480 1 0 $X=316530 $Y=55360
X10304 3 1 DECAP5JI3V $T=316960 60480 0 0 $X=316530 $Y=59840
X10305 3 1 DECAP5JI3V $T=316960 69440 1 0 $X=316530 $Y=64320
X10306 3 1 DECAP5JI3V $T=316960 96320 0 0 $X=316530 $Y=95680
X10307 3 1 DECAP5JI3V $T=316960 105280 1 0 $X=316530 $Y=100160
X10308 3 1 DECAP5JI3V $T=316960 114240 1 0 $X=316530 $Y=109120
X10309 3 1 DECAP5JI3V $T=316960 141120 0 0 $X=316530 $Y=140480
X10310 3 1 DECAP5JI3V $T=316960 150080 0 0 $X=316530 $Y=149440
X10311 3 1 DECAP5JI3V $T=320320 105280 0 0 $X=319890 $Y=104640
X10312 3 1 DECAP5JI3V $T=322000 87360 0 0 $X=321570 $Y=86720
X10313 3 1 DECAP5JI3V $T=322000 114240 0 0 $X=321570 $Y=113600
X10314 3 1 DECAP5JI3V $T=322000 123200 0 0 $X=321570 $Y=122560
X10315 3 1 DECAP5JI3V $T=322000 212800 0 0 $X=321570 $Y=212160
X10316 3 1 DECAP5JI3V $T=323120 132160 0 0 $X=322690 $Y=131520
X10317 3 1 DECAP5JI3V $T=329840 132160 1 180 $X=326610 $Y=131520
X10318 3 1 DECAP5JI3V $T=332080 42560 0 0 $X=331650 $Y=41920
X10319 3 1 DECAP5JI3V $T=333760 132160 0 0 $X=333330 $Y=131520
X10320 3 1 DECAP5JI3V $T=334320 105280 0 0 $X=333890 $Y=104640
X10321 3 1 DECAP5JI3V $T=352800 141120 1 180 $X=349570 $Y=140480
X10322 3 1 DECAP5JI3V $T=357840 132160 0 0 $X=357410 $Y=131520
X10323 3 1 DECAP5JI3V $T=357840 141120 1 0 $X=357410 $Y=136000
X10324 3 1 DECAP5JI3V $T=361200 42560 0 0 $X=360770 $Y=41920
X10325 3 1 DECAP5JI3V $T=361200 51520 1 0 $X=360770 $Y=46400
X10326 3 1 DECAP5JI3V $T=361200 159040 0 0 $X=360770 $Y=158400
X10327 3 1 DECAP5JI3V $T=366240 123200 0 0 $X=365810 $Y=122560
X10328 3 1 DECAP5JI3V $T=422240 24640 0 0 $X=421810 $Y=24000
X10329 3 1 DECAP5JI3V $T=422240 69440 1 0 $X=421810 $Y=64320
X10330 3 1 DECAP5JI3V $T=422240 78400 0 0 $X=421810 $Y=77760
X10331 3 1 DECAP5JI3V $T=422240 87360 0 0 $X=421810 $Y=86720
X10332 3 1 DECAP5JI3V $T=422240 96320 1 0 $X=421810 $Y=91200
X10333 3 1 DECAP5JI3V $T=422240 96320 0 0 $X=421810 $Y=95680
X10334 3 1 DECAP5JI3V $T=422240 105280 1 0 $X=421810 $Y=100160
X10335 3 1 DECAP5JI3V $T=422240 105280 0 0 $X=421810 $Y=104640
X10336 3 1 DECAP5JI3V $T=422240 114240 0 0 $X=421810 $Y=113600
X10337 3 1 DECAP5JI3V $T=422240 123200 1 0 $X=421810 $Y=118080
X10338 3 1 DECAP5JI3V $T=422240 132160 0 0 $X=421810 $Y=131520
X10339 3 1 DECAP5JI3V $T=422240 141120 1 0 $X=421810 $Y=136000
X10340 3 1 DECAP5JI3V $T=422240 150080 0 0 $X=421810 $Y=149440
X10341 3 1 DECAP5JI3V $T=422240 159040 1 0 $X=421810 $Y=153920
X10342 3 1 DECAP5JI3V $T=422240 176960 0 0 $X=421810 $Y=176320
X10343 3 1 DECAP5JI3V $T=422240 185920 1 0 $X=421810 $Y=180800
X10344 3 1 DECAP5JI3V $T=422240 194880 1 0 $X=421810 $Y=189760
X10345 3 1 DECAP5JI3V $T=422240 212800 0 0 $X=421810 $Y=212160
X10346 3 1 DECAP15JI3V $T=20160 33600 1 0 $X=19730 $Y=28480
X10347 3 1 DECAP15JI3V $T=20160 69440 0 0 $X=19730 $Y=68800
X10348 3 1 DECAP15JI3V $T=20160 123200 1 0 $X=19730 $Y=118080
X10349 3 1 DECAP15JI3V $T=20160 194880 1 0 $X=19730 $Y=189760
X10350 3 1 DECAP15JI3V $T=20160 203840 0 0 $X=19730 $Y=203200
X10351 3 1 DECAP15JI3V $T=34160 212800 0 0 $X=33730 $Y=212160
X10352 3 1 DECAP15JI3V $T=70000 33600 0 0 $X=69570 $Y=32960
X10353 3 1 DECAP15JI3V $T=75040 132160 0 0 $X=74610 $Y=131520
X10354 3 1 DECAP15JI3V $T=90720 123200 0 0 $X=90290 $Y=122560
X10355 3 1 DECAP15JI3V $T=100240 150080 0 0 $X=99810 $Y=149440
X10356 3 1 DECAP15JI3V $T=100240 159040 1 0 $X=99810 $Y=153920
X10357 3 1 DECAP15JI3V $T=100800 159040 0 0 $X=100370 $Y=158400
X10358 3 1 DECAP15JI3V $T=104720 114240 0 0 $X=104290 $Y=113600
X10359 3 1 DECAP15JI3V $T=104720 123200 1 0 $X=104290 $Y=118080
X10360 3 1 DECAP15JI3V $T=104720 185920 0 0 $X=104290 $Y=185280
X10361 3 1 DECAP15JI3V $T=104720 194880 1 0 $X=104290 $Y=189760
X10362 3 1 DECAP15JI3V $T=110320 212800 1 0 $X=109890 $Y=207680
X10363 3 1 DECAP15JI3V $T=110320 221760 1 0 $X=109890 $Y=216640
X10364 3 1 DECAP15JI3V $T=134400 87360 1 0 $X=133970 $Y=82240
X10365 3 1 DECAP15JI3V $T=134400 141120 1 0 $X=133970 $Y=136000
X10366 3 1 DECAP15JI3V $T=141120 78400 0 0 $X=140690 $Y=77760
X10367 3 1 DECAP15JI3V $T=148960 114240 1 0 $X=148530 $Y=109120
X10368 3 1 DECAP15JI3V $T=154000 221760 1 0 $X=153570 $Y=216640
X10369 3 1 DECAP15JI3V $T=177520 87360 1 0 $X=177090 $Y=82240
X10370 3 1 DECAP15JI3V $T=186480 78400 0 0 $X=186050 $Y=77760
X10371 3 1 DECAP15JI3V $T=206080 87360 0 0 $X=205650 $Y=86720
X10372 3 1 DECAP15JI3V $T=206080 150080 1 0 $X=205650 $Y=144960
X10373 3 1 DECAP15JI3V $T=206640 141120 1 0 $X=206210 $Y=136000
X10374 3 1 DECAP15JI3V $T=206640 159040 0 0 $X=206210 $Y=158400
X10375 3 1 DECAP15JI3V $T=206640 176960 0 0 $X=206210 $Y=176320
X10376 3 1 DECAP15JI3V $T=207760 96320 1 0 $X=207330 $Y=91200
X10377 3 1 DECAP15JI3V $T=208880 141120 0 0 $X=208450 $Y=140480
X10378 3 1 DECAP15JI3V $T=208880 203840 0 0 $X=208450 $Y=203200
X10379 3 1 DECAP15JI3V $T=210000 203840 1 0 $X=209570 $Y=198720
X10380 3 1 DECAP15JI3V $T=210560 221760 1 0 $X=210130 $Y=216640
X10381 3 1 DECAP15JI3V $T=211120 87360 1 0 $X=210690 $Y=82240
X10382 3 1 DECAP15JI3V $T=259280 96320 1 0 $X=258850 $Y=91200
X10383 3 1 DECAP15JI3V $T=270480 78400 0 0 $X=270050 $Y=77760
X10384 3 1 DECAP15JI3V $T=273840 114240 1 0 $X=273410 $Y=109120
X10385 3 1 DECAP15JI3V $T=279440 150080 0 0 $X=279010 $Y=149440
X10386 3 1 DECAP15JI3V $T=308560 123200 1 0 $X=308130 $Y=118080
X10387 3 1 DECAP15JI3V $T=308560 132160 1 0 $X=308130 $Y=127040
X10388 3 1 DECAP15JI3V $T=309680 87360 0 0 $X=309250 $Y=86720
X10389 3 1 DECAP15JI3V $T=309680 96320 1 0 $X=309250 $Y=91200
X10390 3 1 DECAP15JI3V $T=309680 123200 0 0 $X=309250 $Y=122560
X10391 3 1 DECAP15JI3V $T=311920 105280 0 0 $X=311490 $Y=104640
X10392 3 1 DECAP15JI3V $T=313600 114240 0 0 $X=313170 $Y=113600
X10393 3 1 DECAP15JI3V $T=316400 185920 1 0 $X=315970 $Y=180800
X10394 3 1 DECAP15JI3V $T=316960 51520 1 0 $X=316530 $Y=46400
X10395 3 1 DECAP15JI3V $T=316960 185920 0 0 $X=316530 $Y=185280
X10396 3 1 DECAP15JI3V $T=316960 194880 1 0 $X=316530 $Y=189760
X10397 3 1 DECAP15JI3V $T=332640 221760 1 0 $X=332210 $Y=216640
X10398 3 1 DECAP15JI3V $T=365120 176960 1 0 $X=364690 $Y=171840
X10399 3 1 DECAP15JI3V $T=366240 185920 0 0 $X=365810 $Y=185280
X10400 3 1 DECAP15JI3V $T=378560 78400 1 0 $X=378130 $Y=73280
X10401 3 1 DECAP15JI3V $T=379120 176960 1 0 $X=378690 $Y=171840
X10402 3 1 DECAP15JI3V $T=384720 42560 1 0 $X=384290 $Y=37440
X10403 3 1 DECAP15JI3V $T=384720 42560 0 0 $X=384290 $Y=41920
X10404 3 1 DECAP15JI3V $T=384720 168000 1 0 $X=384290 $Y=162880
X10405 3 1 DECAP15JI3V $T=400960 78400 1 0 $X=400530 $Y=73280
X10406 3 1 DECAP15JI3V $T=400960 87360 1 0 $X=400530 $Y=82240
X10407 3 1 DECAP15JI3V $T=400960 212800 1 0 $X=400530 $Y=207680
X10408 3 1 DECAP15JI3V $T=402080 185920 1 0 $X=401650 $Y=180800
X10409 3 1 DECAP15JI3V $T=404880 203840 0 0 $X=404450 $Y=203200
X10410 3 1 DECAP15JI3V $T=406000 176960 0 0 $X=405570 $Y=176320
X10411 3 1 DECAP15JI3V $T=408800 33600 1 0 $X=408370 $Y=28480
X10412 3 1 DECAP15JI3V $T=408800 114240 1 0 $X=408370 $Y=109120
X10413 3 1 DECAP15JI3V $T=408800 141120 0 0 $X=408370 $Y=140480
X10414 3 1 DECAP15JI3V $T=409920 96320 0 0 $X=409490 $Y=95680
X10415 3 1 DECAP15JI3V $T=409920 105280 1 0 $X=409490 $Y=100160
X10416 3 1 DECAP15JI3V $T=409920 114240 0 0 $X=409490 $Y=113600
X10417 3 1 DECAP15JI3V $T=409920 132160 0 0 $X=409490 $Y=131520
X10418 3 1 DECAP15JI3V $T=409920 141120 1 0 $X=409490 $Y=136000
X10419 3 1 DECAP15JI3V $T=416640 185920 0 0 $X=416210 $Y=185280
D0 2 3 p_ddnwmv AREA=8.4767e-08 PJ=0.00123324 perimeter=0.00123324 $X=17730 $Y=17520 $dt=2
D1 1 3 p_dipdnwmv AREA=1.66597e-09 PJ=0.000831805 perimeter=0.000831805 $X=27180 $Y=94080 $dt=3
D2 1 3 p_dipdnwmv AREA=1.65762e-09 PJ=0.000829452 perimeter=0.000829452 $X=28860 $Y=210560 $dt=3
D3 1 3 p_dipdnwmv AREA=1.66947e-09 PJ=0.000832178 perimeter=0.000832178 $X=40620 $Y=129920 $dt=3
D4 1 3 p_dipdnwmv AREA=1.65893e-09 PJ=0.000835699 perimeter=0.000835699 $X=53650 $Y=174710 $dt=3
D5 1 3 p_dipdnwmv AREA=1.6774e-09 PJ=0.000833895 perimeter=0.000833895 $X=57010 $Y=67190 $dt=3
D6 1 3 p_dipdnwmv AREA=1.62356e-09 PJ=0.000824013 perimeter=0.000824013 $X=91990 $Y=192430 $dt=3
D7 1 3 p_dipdnwmv AREA=1.66696e-09 PJ=0.000835085 perimeter=0.000835085 $X=101900 $Y=85110 $dt=3
D8 1 3 p_dipdnwmv AREA=1.65811e-09 PJ=0.000830245 perimeter=0.000830245 $X=101900 $Y=103030 $dt=3
D9 1 3 p_dipdnwmv AREA=1.66166e-09 PJ=0.000833269 perimeter=0.000833269 $X=101900 $Y=147830 $dt=3
D10 1 3 p_dipdnwmv AREA=1.6681e-09 PJ=0.000833335 perimeter=0.000833335 $X=113570 $Y=76150 $dt=3
D11 1 3 p_dipdnwmv AREA=1.66771e-09 PJ=0.000832586 perimeter=0.000832586 $X=118050 $Y=120950 $dt=3
D12 1 3 p_dipdnwmv AREA=1.6716e-09 PJ=0.000833709 perimeter=0.000833709 $X=143250 $Y=138870 $dt=3
D13 1 3 p_dipdnwmv AREA=1.66525e-09 PJ=0.000831652 perimeter=0.000831652 $X=143810 $Y=111990 $dt=3
D14 1 3 p_dipdnwmv AREA=1.67857e-09 PJ=0.000836374 perimeter=0.000836374 $X=144370 $Y=49270 $dt=3
D15 1 3 p_dipdnwmv AREA=1.67238e-09 PJ=0.000835208 perimeter=0.000835208 $X=146050 $Y=165750 $dt=3
D16 1 3 p_dipdnwmv AREA=1.66036e-09 PJ=0.000835202 perimeter=0.000835202 $X=161170 $Y=40310 $dt=3
D17 1 3 p_dipdnwmv AREA=1.67755e-09 PJ=0.000834786 perimeter=0.000834786 $X=164530 $Y=156790 $dt=3
D18 1 3 p_dipdnwmv AREA=1.08218e-09 PJ=0.000821773 perimeter=0.000821773 $X=164530 $Y=219510 $dt=3
D19 1 3 p_dipdnwmv AREA=1.6798e-09 PJ=0.000840932 perimeter=0.000840932 $X=179090 $Y=58230 $dt=3
D20 1 3 p_dipdnwmv AREA=1.6264e-09 PJ=0.000826294 perimeter=0.000826294 $X=189730 $Y=31350 $dt=3
D21 1 3 p_dipdnwmv AREA=1.6322e-09 PJ=0.00082472 perimeter=0.00082472 $X=207740 $Y=183670 $dt=3
D22 1 3 p_dipdnwmv AREA=1.61051e-09 PJ=0.000822069 perimeter=0.000822069 $X=273360 $Y=22480 $dt=3
D23 1 3 p_dipdnwmv AREA=1.63119e-09 PJ=0.000824905 perimeter=0.000824905 $X=273880 $Y=201390 $dt=3
.ends aska_dig
